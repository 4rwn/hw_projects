module sorter #(
    parameter VALUE_BITS = 8,
    parameter DEPTH = 5,
    parameter DIRECTION = 0,
    parameter SIZE = 1 << DEPTH // Do not override
) (
    input logic clk,

    input logic [SIZE-1:0][VALUE_BITS-1:0] in,
    output logic [SIZE-1:0][VALUE_BITS-1:0] out
);
    genvar i;
    generate
        if (DEPTH > 5) begin
            logic [SIZE-1:0][VALUE_BITS-1:0] intermediate;

            sorter #(
                .VALUE_BITS(VALUE_BITS),
                .DEPTH(DEPTH - 1),
                .DIRECTION(DIRECTION)
            ) first_sorter (
                .clk(clk),

                .in(in[SIZE/2-1:0]),
                .out(intermediate[SIZE/2-1:0])
            );

            sorter #(
                .VALUE_BITS(VALUE_BITS),
                .DEPTH(DEPTH - 1),
                .DIRECTION(1 - DIRECTION)
            ) second_sorter (
                .clk(clk),
                
                .in(in[SIZE-1:SIZE/2]),
                .out(intermediate[SIZE-1:SIZE/2])
            );

            merger #(
                .VALUE_BITS(VALUE_BITS),
                .DEPTH(DEPTH),
                .DIRECTION(DIRECTION)
            ) merger (
                .clk(clk),

                .in(intermediate),
                .out(out)
            );
        end else begin
            logic [31:0][VALUE_BITS-1:0] t0;
            logic [31:0][VALUE_BITS-1:0] t1;
            logic [31:0][VALUE_BITS-1:0] t2;
            logic [31:0][VALUE_BITS-1:0] t3;
            logic [31:0][VALUE_BITS-1:0] t4;
            logic [31:0][VALUE_BITS-1:0] t5;
            logic [31:0][VALUE_BITS-1:0] t6;
            logic [31:0][VALUE_BITS-1:0] t7;
            logic [31:0][VALUE_BITS-1:0] t8;
            logic [31:0][VALUE_BITS-1:0] t9;
            logic [31:0][VALUE_BITS-1:0] t10;
            logic [31:0][VALUE_BITS-1:0] t11;
            logic [31:0][VALUE_BITS-1:0] t12;
            logic [31:0][VALUE_BITS-1:0] t13;
            assign {t0[0], t0[1]} = (in[0] > in[1]) ? {in[1], in[0]} : {in[0], in[1]};
            assign {t0[2], t0[3]} = (in[2] > in[3]) ? {in[3], in[2]} : {in[2], in[3]};
            assign {t0[4], t0[5]} = (in[4] > in[5]) ? {in[5], in[4]} : {in[4], in[5]};
            assign {t0[6], t0[7]} = (in[6] > in[7]) ? {in[7], in[6]} : {in[6], in[7]};
            assign {t0[8], t0[9]} = (in[8] > in[9]) ? {in[9], in[8]} : {in[8], in[9]};
            assign {t0[10], t0[11]} = (in[10] > in[11]) ? {in[11], in[10]} : {in[10], in[11]};
            assign {t0[12], t0[13]} = (in[12] > in[13]) ? {in[13], in[12]} : {in[12], in[13]};
            assign {t0[14], t0[15]} = (in[14] > in[15]) ? {in[15], in[14]} : {in[14], in[15]};
            assign {t0[16], t0[17]} = (in[16] > in[17]) ? {in[17], in[16]} : {in[16], in[17]};
            assign {t0[18], t0[19]} = (in[18] > in[19]) ? {in[19], in[18]} : {in[18], in[19]};
            assign {t0[20], t0[21]} = (in[20] > in[21]) ? {in[21], in[20]} : {in[20], in[21]};
            assign {t0[22], t0[23]} = (in[22] > in[23]) ? {in[23], in[22]} : {in[22], in[23]};
            assign {t0[24], t0[25]} = (in[24] > in[25]) ? {in[25], in[24]} : {in[24], in[25]};
            assign {t0[26], t0[27]} = (in[26] > in[27]) ? {in[27], in[26]} : {in[26], in[27]};
            assign {t0[28], t0[29]} = (in[28] > in[29]) ? {in[29], in[28]} : {in[28], in[29]};
            assign {t0[30], t0[31]} = (in[30] > in[31]) ? {in[31], in[30]} : {in[30], in[31]};
            assign {t1[0], t1[2]} = (t0[0] > t0[2]) ? {t0[2], t0[0]} : {t0[0], t0[2]};
            assign {t1[1], t1[3]} = (t0[1] > t0[3]) ? {t0[3], t0[1]} : {t0[1], t0[3]};
            assign {t1[4], t1[6]} = (t0[4] > t0[6]) ? {t0[6], t0[4]} : {t0[4], t0[6]};
            assign {t1[5], t1[7]} = (t0[5] > t0[7]) ? {t0[7], t0[5]} : {t0[5], t0[7]};
            assign {t1[8], t1[10]} = (t0[8] > t0[10]) ? {t0[10], t0[8]} : {t0[8], t0[10]};
            assign {t1[9], t1[11]} = (t0[9] > t0[11]) ? {t0[11], t0[9]} : {t0[9], t0[11]};
            assign {t1[12], t1[14]} = (t0[12] > t0[14]) ? {t0[14], t0[12]} : {t0[12], t0[14]};
            assign {t1[13], t1[15]} = (t0[13] > t0[15]) ? {t0[15], t0[13]} : {t0[13], t0[15]};
            assign {t1[16], t1[18]} = (t0[16] > t0[18]) ? {t0[18], t0[16]} : {t0[16], t0[18]};
            assign {t1[17], t1[19]} = (t0[17] > t0[19]) ? {t0[19], t0[17]} : {t0[17], t0[19]};
            assign {t1[20], t1[22]} = (t0[20] > t0[22]) ? {t0[22], t0[20]} : {t0[20], t0[22]};
            assign {t1[21], t1[23]} = (t0[21] > t0[23]) ? {t0[23], t0[21]} : {t0[21], t0[23]};
            assign {t1[24], t1[26]} = (t0[24] > t0[26]) ? {t0[26], t0[24]} : {t0[24], t0[26]};
            assign {t1[25], t1[27]} = (t0[25] > t0[27]) ? {t0[27], t0[25]} : {t0[25], t0[27]};
            assign {t1[28], t1[30]} = (t0[28] > t0[30]) ? {t0[30], t0[28]} : {t0[28], t0[30]};
            assign {t1[29], t1[31]} = (t0[29] > t0[31]) ? {t0[31], t0[29]} : {t0[29], t0[31]};
            assign {t2[0], t2[4]} = (t1[0] > t1[4]) ? {t1[4], t1[0]} : {t1[0], t1[4]};
            assign {t2[1], t2[5]} = (t1[1] > t1[5]) ? {t1[5], t1[1]} : {t1[1], t1[5]};
            assign {t2[2], t2[6]} = (t1[2] > t1[6]) ? {t1[6], t1[2]} : {t1[2], t1[6]};
            assign {t2[3], t2[7]} = (t1[3] > t1[7]) ? {t1[7], t1[3]} : {t1[3], t1[7]};
            assign {t2[8], t2[12]} = (t1[8] > t1[12]) ? {t1[12], t1[8]} : {t1[8], t1[12]};
            assign {t2[9], t2[13]} = (t1[9] > t1[13]) ? {t1[13], t1[9]} : {t1[9], t1[13]};
            assign {t2[10], t2[14]} = (t1[10] > t1[14]) ? {t1[14], t1[10]} : {t1[10], t1[14]};
            assign {t2[11], t2[15]} = (t1[11] > t1[15]) ? {t1[15], t1[11]} : {t1[11], t1[15]};
            assign {t2[16], t2[20]} = (t1[16] > t1[20]) ? {t1[20], t1[16]} : {t1[16], t1[20]};
            assign {t2[17], t2[21]} = (t1[17] > t1[21]) ? {t1[21], t1[17]} : {t1[17], t1[21]};
            assign {t2[18], t2[22]} = (t1[18] > t1[22]) ? {t1[22], t1[18]} : {t1[18], t1[22]};
            assign {t2[19], t2[23]} = (t1[19] > t1[23]) ? {t1[23], t1[19]} : {t1[19], t1[23]};
            assign {t2[24], t2[28]} = (t1[24] > t1[28]) ? {t1[28], t1[24]} : {t1[24], t1[28]};
            assign {t2[25], t2[29]} = (t1[25] > t1[29]) ? {t1[29], t1[25]} : {t1[25], t1[29]};
            assign {t2[26], t2[30]} = (t1[26] > t1[30]) ? {t1[30], t1[26]} : {t1[26], t1[30]};
            assign {t2[27], t2[31]} = (t1[27] > t1[31]) ? {t1[31], t1[27]} : {t1[27], t1[31]};
            assign {t3[0], t3[8]} = (t2[0] > t2[8]) ? {t2[8], t2[0]} : {t2[0], t2[8]};
            assign {t3[1], t3[9]} = (t2[1] > t2[9]) ? {t2[9], t2[1]} : {t2[1], t2[9]};
            assign {t3[2], t3[10]} = (t2[2] > t2[10]) ? {t2[10], t2[2]} : {t2[2], t2[10]};
            assign {t3[3], t3[11]} = (t2[3] > t2[11]) ? {t2[11], t2[3]} : {t2[3], t2[11]};
            assign {t3[4], t3[12]} = (t2[4] > t2[12]) ? {t2[12], t2[4]} : {t2[4], t2[12]};
            assign {t3[5], t3[13]} = (t2[5] > t2[13]) ? {t2[13], t2[5]} : {t2[5], t2[13]};
            assign {t3[6], t3[14]} = (t2[6] > t2[14]) ? {t2[14], t2[6]} : {t2[6], t2[14]};
            assign {t3[7], t3[15]} = (t2[7] > t2[15]) ? {t2[15], t2[7]} : {t2[7], t2[15]};
            assign {t3[16], t3[24]} = (t2[16] > t2[24]) ? {t2[24], t2[16]} : {t2[16], t2[24]};
            assign {t3[17], t3[25]} = (t2[17] > t2[25]) ? {t2[25], t2[17]} : {t2[17], t2[25]};
            assign {t3[18], t3[26]} = (t2[18] > t2[26]) ? {t2[26], t2[18]} : {t2[18], t2[26]};
            assign {t3[19], t3[27]} = (t2[19] > t2[27]) ? {t2[27], t2[19]} : {t2[19], t2[27]};
            assign {t3[20], t3[28]} = (t2[20] > t2[28]) ? {t2[28], t2[20]} : {t2[20], t2[28]};
            assign {t3[21], t3[29]} = (t2[21] > t2[29]) ? {t2[29], t2[21]} : {t2[21], t2[29]};
            assign {t3[22], t3[30]} = (t2[22] > t2[30]) ? {t2[30], t2[22]} : {t2[22], t2[30]};
            assign {t3[23], t3[31]} = (t2[23] > t2[31]) ? {t2[31], t2[23]} : {t2[23], t2[31]};
            assign {t4[0], t4[16]} = (t3[0] > t3[16]) ? {t3[16], t3[0]} : {t3[0], t3[16]};
            assign {t4[1], t4[8]} = (t3[1] > t3[8]) ? {t3[8], t3[1]} : {t3[1], t3[8]};
            assign {t4[2], t4[4]} = (t3[2] > t3[4]) ? {t3[4], t3[2]} : {t3[2], t3[4]};
            assign {t4[3], t4[12]} = (t3[3] > t3[12]) ? {t3[12], t3[3]} : {t3[3], t3[12]};
            assign {t4[5], t4[10]} = (t3[5] > t3[10]) ? {t3[10], t3[5]} : {t3[5], t3[10]};
            assign {t4[6], t4[9]} = (t3[6] > t3[9]) ? {t3[9], t3[6]} : {t3[6], t3[9]};
            assign {t4[7], t4[14]} = (t3[7] > t3[14]) ? {t3[14], t3[7]} : {t3[7], t3[14]};
            assign {t4[11], t4[13]} = (t3[11] > t3[13]) ? {t3[13], t3[11]} : {t3[11], t3[13]};
            assign {t4[15], t4[31]} = (t3[15] > t3[31]) ? {t3[31], t3[15]} : {t3[15], t3[31]};
            assign {t4[17], t4[24]} = (t3[17] > t3[24]) ? {t3[24], t3[17]} : {t3[17], t3[24]};
            assign {t4[18], t4[20]} = (t3[18] > t3[20]) ? {t3[20], t3[18]} : {t3[18], t3[20]};
            assign {t4[19], t4[28]} = (t3[19] > t3[28]) ? {t3[28], t3[19]} : {t3[19], t3[28]};
            assign {t4[21], t4[26]} = (t3[21] > t3[26]) ? {t3[26], t3[21]} : {t3[21], t3[26]};
            assign {t4[22], t4[25]} = (t3[22] > t3[25]) ? {t3[25], t3[22]} : {t3[22], t3[25]};
            assign {t4[23], t4[30]} = (t3[23] > t3[30]) ? {t3[30], t3[23]} : {t3[23], t3[30]};
            assign {t4[27], t4[29]} = (t3[27] > t3[29]) ? {t3[29], t3[27]} : {t3[27], t3[29]};
            assign {t5[1], t5[2]} = (t4[1] > t4[2]) ? {t4[2], t4[1]} : {t4[1], t4[2]};
            assign {t5[3], t5[5]} = (t4[3] > t4[5]) ? {t4[5], t4[3]} : {t4[3], t4[5]};
            assign {t5[4], t5[8]} = (t4[4] > t4[8]) ? {t4[8], t4[4]} : {t4[4], t4[8]};
            assign {t5[6], t5[22]} = (t4[6] > t4[22]) ? {t4[22], t4[6]} : {t4[6], t4[22]};
            assign {t5[7], t5[11]} = (t4[7] > t4[11]) ? {t4[11], t4[7]} : {t4[7], t4[11]};
            assign {t5[9], t5[25]} = (t4[9] > t4[25]) ? {t4[25], t4[9]} : {t4[9], t4[25]};
            assign {t5[10], t5[12]} = (t4[10] > t4[12]) ? {t4[12], t4[10]} : {t4[10], t4[12]};
            assign {t5[13], t5[14]} = (t4[13] > t4[14]) ? {t4[14], t4[13]} : {t4[13], t4[14]};
            assign {t5[17], t5[18]} = (t4[17] > t4[18]) ? {t4[18], t4[17]} : {t4[17], t4[18]};
            assign {t5[19], t5[21]} = (t4[19] > t4[21]) ? {t4[21], t4[19]} : {t4[19], t4[21]};
            assign {t5[20], t5[24]} = (t4[20] > t4[24]) ? {t4[24], t4[20]} : {t4[20], t4[24]};
            assign {t5[23], t5[27]} = (t4[23] > t4[27]) ? {t4[27], t4[23]} : {t4[23], t4[27]};
            assign {t5[26], t5[28]} = (t4[26] > t4[28]) ? {t4[28], t4[26]} : {t4[26], t4[28]};
            assign {t5[29], t5[30]} = (t4[29] > t4[30]) ? {t4[30], t4[29]} : {t4[29], t4[30]};
            assign t5[0] = t4[0];
            assign t5[15] = t4[15];
            assign t5[16] = t4[16];
            assign t5[31] = t4[31];
            assign {t6[1], t6[17]} = (t5[1] > t5[17]) ? {t5[17], t5[1]} : {t5[1], t5[17]};
            assign {t6[2], t6[18]} = (t5[2] > t5[18]) ? {t5[18], t5[2]} : {t5[2], t5[18]};
            assign {t6[3], t6[19]} = (t5[3] > t5[19]) ? {t5[19], t5[3]} : {t5[3], t5[19]};
            assign {t6[4], t6[20]} = (t5[4] > t5[20]) ? {t5[20], t5[4]} : {t5[4], t5[20]};
            assign {t6[5], t6[10]} = (t5[5] > t5[10]) ? {t5[10], t5[5]} : {t5[5], t5[10]};
            assign {t6[7], t6[23]} = (t5[7] > t5[23]) ? {t5[23], t5[7]} : {t5[7], t5[23]};
            assign {t6[8], t6[24]} = (t5[8] > t5[24]) ? {t5[24], t5[8]} : {t5[8], t5[24]};
            assign {t6[11], t6[27]} = (t5[11] > t5[27]) ? {t5[27], t5[11]} : {t5[11], t5[27]};
            assign {t6[12], t6[28]} = (t5[12] > t5[28]) ? {t5[28], t5[12]} : {t5[12], t5[28]};
            assign {t6[13], t6[29]} = (t5[13] > t5[29]) ? {t5[29], t5[13]} : {t5[13], t5[29]};
            assign {t6[14], t6[30]} = (t5[14] > t5[30]) ? {t5[30], t5[14]} : {t5[14], t5[30]};
            assign {t6[21], t6[26]} = (t5[21] > t5[26]) ? {t5[26], t5[21]} : {t5[21], t5[26]};
            assign t6[0] = t5[0];
            assign t6[6] = t5[6];
            assign t6[9] = t5[9];
            assign t6[15] = t5[15];
            assign t6[16] = t5[16];
            assign t6[22] = t5[22];
            assign t6[25] = t5[25];
            assign t6[31] = t5[31];
            assign {t7[3], t7[17]} = (t6[3] > t6[17]) ? {t6[17], t6[3]} : {t6[3], t6[17]};
            assign {t7[4], t7[16]} = (t6[4] > t6[16]) ? {t6[16], t6[4]} : {t6[4], t6[16]};
            assign {t7[5], t7[21]} = (t6[5] > t6[21]) ? {t6[21], t6[5]} : {t6[5], t6[21]};
            assign {t7[6], t7[18]} = (t6[6] > t6[18]) ? {t6[18], t6[6]} : {t6[6], t6[18]};
            assign {t7[7], t7[9]} = (t6[7] > t6[9]) ? {t6[9], t6[7]} : {t6[7], t6[9]};
            assign {t7[8], t7[20]} = (t6[8] > t6[20]) ? {t6[20], t6[8]} : {t6[8], t6[20]};
            assign {t7[10], t7[26]} = (t6[10] > t6[26]) ? {t6[26], t6[10]} : {t6[10], t6[26]};
            assign {t7[11], t7[23]} = (t6[11] > t6[23]) ? {t6[23], t6[11]} : {t6[11], t6[23]};
            assign {t7[13], t7[25]} = (t6[13] > t6[25]) ? {t6[25], t6[13]} : {t6[13], t6[25]};
            assign {t7[14], t7[28]} = (t6[14] > t6[28]) ? {t6[28], t6[14]} : {t6[14], t6[28]};
            assign {t7[15], t7[27]} = (t6[15] > t6[27]) ? {t6[27], t6[15]} : {t6[15], t6[27]};
            assign {t7[22], t7[24]} = (t6[22] > t6[24]) ? {t6[24], t6[22]} : {t6[22], t6[24]};
            assign t7[0] = t6[0];
            assign t7[1] = t6[1];
            assign t7[2] = t6[2];
            assign t7[12] = t6[12];
            assign t7[19] = t6[19];
            assign t7[29] = t6[29];
            assign t7[30] = t6[30];
            assign t7[31] = t6[31];
            assign {t8[1], t8[4]} = (t7[1] > t7[4]) ? {t7[4], t7[1]} : {t7[1], t7[4]};
            assign {t8[3], t8[8]} = (t7[3] > t7[8]) ? {t7[8], t7[3]} : {t7[3], t7[8]};
            assign {t8[5], t8[16]} = (t7[5] > t7[16]) ? {t7[16], t7[5]} : {t7[5], t7[16]};
            assign {t8[7], t8[17]} = (t7[7] > t7[17]) ? {t7[17], t7[7]} : {t7[7], t7[17]};
            assign {t8[9], t8[21]} = (t7[9] > t7[21]) ? {t7[21], t7[9]} : {t7[9], t7[21]};
            assign {t8[10], t8[22]} = (t7[10] > t7[22]) ? {t7[22], t7[10]} : {t7[10], t7[22]};
            assign {t8[11], t8[19]} = (t7[11] > t7[19]) ? {t7[19], t7[11]} : {t7[11], t7[19]};
            assign {t8[12], t8[20]} = (t7[12] > t7[20]) ? {t7[20], t7[12]} : {t7[12], t7[20]};
            assign {t8[14], t8[24]} = (t7[14] > t7[24]) ? {t7[24], t7[14]} : {t7[14], t7[24]};
            assign {t8[15], t8[26]} = (t7[15] > t7[26]) ? {t7[26], t7[15]} : {t7[15], t7[26]};
            assign {t8[23], t8[28]} = (t7[23] > t7[28]) ? {t7[28], t7[23]} : {t7[23], t7[28]};
            assign {t8[27], t8[30]} = (t7[27] > t7[30]) ? {t7[30], t7[27]} : {t7[27], t7[30]};
            assign t8[0] = t7[0];
            assign t8[2] = t7[2];
            assign t8[6] = t7[6];
            assign t8[13] = t7[13];
            assign t8[18] = t7[18];
            assign t8[25] = t7[25];
            assign t8[29] = t7[29];
            assign t8[31] = t7[31];
            assign {t9[2], t9[5]} = (t8[2] > t8[5]) ? {t8[5], t8[2]} : {t8[2], t8[5]};
            assign {t9[7], t9[8]} = (t8[7] > t8[8]) ? {t8[8], t8[7]} : {t8[7], t8[8]};
            assign {t9[9], t9[18]} = (t8[9] > t8[18]) ? {t8[18], t8[9]} : {t8[9], t8[18]};
            assign {t9[11], t9[17]} = (t8[11] > t8[17]) ? {t8[17], t8[11]} : {t8[11], t8[17]};
            assign {t9[12], t9[16]} = (t8[12] > t8[16]) ? {t8[16], t8[12]} : {t8[12], t8[16]};
            assign {t9[13], t9[22]} = (t8[13] > t8[22]) ? {t8[22], t8[13]} : {t8[13], t8[22]};
            assign {t9[14], t9[20]} = (t8[14] > t8[20]) ? {t8[20], t8[14]} : {t8[14], t8[20]};
            assign {t9[15], t9[19]} = (t8[15] > t8[19]) ? {t8[19], t8[15]} : {t8[15], t8[19]};
            assign {t9[23], t9[24]} = (t8[23] > t8[24]) ? {t8[24], t8[23]} : {t8[23], t8[24]};
            assign {t9[26], t9[29]} = (t8[26] > t8[29]) ? {t8[29], t8[26]} : {t8[26], t8[29]};
            assign t9[0] = t8[0];
            assign t9[1] = t8[1];
            assign t9[3] = t8[3];
            assign t9[4] = t8[4];
            assign t9[6] = t8[6];
            assign t9[10] = t8[10];
            assign t9[21] = t8[21];
            assign t9[25] = t8[25];
            assign t9[27] = t8[27];
            assign t9[28] = t8[28];
            assign t9[30] = t8[30];
            assign t9[31] = t8[31];
            assign {t10[2], t10[4]} = (t9[2] > t9[4]) ? {t9[4], t9[2]} : {t9[2], t9[4]};
            assign {t10[6], t10[12]} = (t9[6] > t9[12]) ? {t9[12], t9[6]} : {t9[6], t9[12]};
            assign {t10[9], t10[16]} = (t9[9] > t9[16]) ? {t9[16], t9[9]} : {t9[9], t9[16]};
            assign {t10[10], t10[11]} = (t9[10] > t9[11]) ? {t9[11], t9[10]} : {t9[10], t9[11]};
            assign {t10[13], t10[17]} = (t9[13] > t9[17]) ? {t9[17], t9[13]} : {t9[13], t9[17]};
            assign {t10[14], t10[18]} = (t9[14] > t9[18]) ? {t9[18], t9[14]} : {t9[14], t9[18]};
            assign {t10[15], t10[22]} = (t9[15] > t9[22]) ? {t9[22], t9[15]} : {t9[15], t9[22]};
            assign {t10[19], t10[25]} = (t9[19] > t9[25]) ? {t9[25], t9[19]} : {t9[19], t9[25]};
            assign {t10[20], t10[21]} = (t9[20] > t9[21]) ? {t9[21], t9[20]} : {t9[20], t9[21]};
            assign {t10[27], t10[29]} = (t9[27] > t9[29]) ? {t9[29], t9[27]} : {t9[27], t9[29]};
            assign t10[0] = t9[0];
            assign t10[1] = t9[1];
            assign t10[3] = t9[3];
            assign t10[5] = t9[5];
            assign t10[7] = t9[7];
            assign t10[8] = t9[8];
            assign t10[23] = t9[23];
            assign t10[24] = t9[24];
            assign t10[26] = t9[26];
            assign t10[28] = t9[28];
            assign t10[30] = t9[30];
            assign t10[31] = t9[31];
            assign {t11[5], t11[6]} = (t10[5] > t10[6]) ? {t10[6], t10[5]} : {t10[5], t10[6]};
            assign {t11[8], t11[12]} = (t10[8] > t10[12]) ? {t10[12], t10[8]} : {t10[8], t10[12]};
            assign {t11[9], t11[10]} = (t10[9] > t10[10]) ? {t10[10], t10[9]} : {t10[9], t10[10]};
            assign {t11[11], t11[13]} = (t10[11] > t10[13]) ? {t10[13], t10[11]} : {t10[11], t10[13]};
            assign {t11[14], t11[16]} = (t10[14] > t10[16]) ? {t10[16], t10[14]} : {t10[14], t10[16]};
            assign {t11[15], t11[17]} = (t10[15] > t10[17]) ? {t10[17], t10[15]} : {t10[15], t10[17]};
            assign {t11[18], t11[20]} = (t10[18] > t10[20]) ? {t10[20], t10[18]} : {t10[18], t10[20]};
            assign {t11[19], t11[23]} = (t10[19] > t10[23]) ? {t10[23], t10[19]} : {t10[19], t10[23]};
            assign {t11[21], t11[22]} = (t10[21] > t10[22]) ? {t10[22], t10[21]} : {t10[21], t10[22]};
            assign {t11[25], t11[26]} = (t10[25] > t10[26]) ? {t10[26], t10[25]} : {t10[25], t10[26]};
            assign t11[0] = t10[0];
            assign t11[1] = t10[1];
            assign t11[2] = t10[2];
            assign t11[3] = t10[3];
            assign t11[4] = t10[4];
            assign t11[7] = t10[7];
            assign t11[24] = t10[24];
            assign t11[27] = t10[27];
            assign t11[28] = t10[28];
            assign t11[29] = t10[29];
            assign t11[30] = t10[30];
            assign t11[31] = t10[31];
            assign {t12[3], t12[5]} = (t11[3] > t11[5]) ? {t11[5], t11[3]} : {t11[3], t11[5]};
            assign {t12[6], t12[7]} = (t11[6] > t11[7]) ? {t11[7], t11[6]} : {t11[6], t11[7]};
            assign {t12[8], t12[9]} = (t11[8] > t11[9]) ? {t11[9], t11[8]} : {t11[8], t11[9]};
            assign {t12[10], t12[12]} = (t11[10] > t11[12]) ? {t11[12], t11[10]} : {t11[10], t11[12]};
            assign {t12[11], t12[14]} = (t11[11] > t11[14]) ? {t11[14], t11[11]} : {t11[11], t11[14]};
            assign {t12[13], t12[16]} = (t11[13] > t11[16]) ? {t11[16], t11[13]} : {t11[13], t11[16]};
            assign {t12[15], t12[18]} = (t11[15] > t11[18]) ? {t11[18], t11[15]} : {t11[15], t11[18]};
            assign {t12[17], t12[20]} = (t11[17] > t11[20]) ? {t11[20], t11[17]} : {t11[17], t11[20]};
            assign {t12[19], t12[21]} = (t11[19] > t11[21]) ? {t11[21], t11[19]} : {t11[19], t11[21]};
            assign {t12[22], t12[23]} = (t11[22] > t11[23]) ? {t11[23], t11[22]} : {t11[22], t11[23]};
            assign {t12[24], t12[25]} = (t11[24] > t11[25]) ? {t11[25], t11[24]} : {t11[24], t11[25]};
            assign {t12[26], t12[28]} = (t11[26] > t11[28]) ? {t11[28], t11[26]} : {t11[26], t11[28]};
            assign t12[0] = t11[0];
            assign t12[1] = t11[1];
            assign t12[2] = t11[2];
            assign t12[4] = t11[4];
            assign t12[27] = t11[27];
            assign t12[29] = t11[29];
            assign t12[30] = t11[30];
            assign t12[31] = t11[31];
            assign {t13[3], t13[4]} = (t12[3] > t12[4]) ? {t12[4], t12[3]} : {t12[3], t12[4]};
            assign {t13[5], t13[6]} = (t12[5] > t12[6]) ? {t12[6], t12[5]} : {t12[5], t12[6]};
            assign {t13[7], t13[8]} = (t12[7] > t12[8]) ? {t12[8], t12[7]} : {t12[7], t12[8]};
            assign {t13[9], t13[10]} = (t12[9] > t12[10]) ? {t12[10], t12[9]} : {t12[9], t12[10]};
            assign {t13[11], t13[12]} = (t12[11] > t12[12]) ? {t12[12], t12[11]} : {t12[11], t12[12]};
            assign {t13[13], t13[14]} = (t12[13] > t12[14]) ? {t12[14], t12[13]} : {t12[13], t12[14]};
            assign {t13[15], t13[16]} = (t12[15] > t12[16]) ? {t12[16], t12[15]} : {t12[15], t12[16]};
            assign {t13[17], t13[18]} = (t12[17] > t12[18]) ? {t12[18], t12[17]} : {t12[17], t12[18]};
            assign {t13[19], t13[20]} = (t12[19] > t12[20]) ? {t12[20], t12[19]} : {t12[19], t12[20]};
            assign {t13[21], t13[22]} = (t12[21] > t12[22]) ? {t12[22], t12[21]} : {t12[21], t12[22]};
            assign {t13[23], t13[24]} = (t12[23] > t12[24]) ? {t12[24], t12[23]} : {t12[23], t12[24]};
            assign {t13[25], t13[26]} = (t12[25] > t12[26]) ? {t12[26], t12[25]} : {t12[25], t12[26]};
            assign {t13[27], t13[28]} = (t12[27] > t12[28]) ? {t12[28], t12[27]} : {t12[27], t12[28]};
            assign t13[0] = t12[0];
            assign t13[1] = t12[1];
            assign t13[2] = t12[2];
            assign t13[29] = t12[29];
            assign t13[30] = t12[30];
            assign t13[31] = t12[31];

            if (DIRECTION == 0) begin
                always_ff @( posedge clk ) begin
                    out <= t13;
                end 
            end else begin
                for (i = 0; i < SIZE; i++) begin
                    always_ff @ ( posedge clk ) begin
                        out[i] <= t13[SIZE-i-1];
                    end
                end
            end
        end
    endgenerate
endmodule