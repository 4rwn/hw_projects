module sorter #(
    parameter VALUE_BITS = 8,
    parameter DEPTH = 6,
    parameter DIRECTION = 0,
    parameter SIZE = 1 << DEPTH // Do not override
) (
    input logic clk,

    input logic [SIZE-1:0][VALUE_BITS-1:0] in,
    output logic [SIZE-1:0][VALUE_BITS-1:0] out
);
    genvar i;
    generate
        if (DEPTH > 6) begin
            logic [SIZE-1:0][VALUE_BITS-1:0] intermediate;

            sorter #(
                .VALUE_BITS(VALUE_BITS),
                .DEPTH(DEPTH - 1),
                .DIRECTION(DIRECTION)
            ) first_sorter (
                .clk(clk),

                .in(in[SIZE/2-1:0]),
                .out(intermediate[SIZE/2-1:0])
            );

            sorter #(
                .VALUE_BITS(VALUE_BITS),
                .DEPTH(DEPTH - 1),
                .DIRECTION(1 - DIRECTION)
            ) second_sorter (
                .clk(clk),
                
                .in(in[SIZE-1:SIZE/2]),
                .out(intermediate[SIZE-1:SIZE/2])
            );

            merger #(
                .VALUE_BITS(VALUE_BITS),
                .DEPTH(DEPTH),
                .DIRECTION(DIRECTION)
            ) merger (
                .clk(clk),

                .in(intermediate),
                .out(out)
            );
        end else begin
            logic [63:0][VALUE_BITS-1:0] t0;
            logic [63:0][VALUE_BITS-1:0] t1;
            logic [63:0][VALUE_BITS-1:0] t2;
            logic [63:0][VALUE_BITS-1:0] t3;
            logic [63:0][VALUE_BITS-1:0] t4;
            logic [63:0][VALUE_BITS-1:0] t5;
            logic [63:0][VALUE_BITS-1:0] t6;
            logic [63:0][VALUE_BITS-1:0] t7;
            logic [63:0][VALUE_BITS-1:0] t8;
            logic [63:0][VALUE_BITS-1:0] t9;
            logic [63:0][VALUE_BITS-1:0] t10;
            logic [63:0][VALUE_BITS-1:0] t11;
            logic [63:0][VALUE_BITS-1:0] t12;
            logic [63:0][VALUE_BITS-1:0] t13;
            logic [63:0][VALUE_BITS-1:0] t14;
            logic [63:0][VALUE_BITS-1:0] t15;
            logic [63:0][VALUE_BITS-1:0] t16;
            logic [63:0][VALUE_BITS-1:0] t17;
            logic [63:0][VALUE_BITS-1:0] t18;
            logic [63:0][VALUE_BITS-1:0] t19;
            assign {t0[0], t0[2]} = (in[0] > in[2]) ? {in[2], in[0]} : {in[0], in[2]};
            assign {t0[1], t0[3]} = (in[1] > in[3]) ? {in[3], in[1]} : {in[1], in[3]};
            assign {t0[4], t0[6]} = (in[4] > in[6]) ? {in[6], in[4]} : {in[4], in[6]};
            assign {t0[5], t0[7]} = (in[5] > in[7]) ? {in[7], in[5]} : {in[5], in[7]};
            assign {t0[8], t0[10]} = (in[8] > in[10]) ? {in[10], in[8]} : {in[8], in[10]};
            assign {t0[9], t0[11]} = (in[9] > in[11]) ? {in[11], in[9]} : {in[9], in[11]};
            assign {t0[12], t0[14]} = (in[12] > in[14]) ? {in[14], in[12]} : {in[12], in[14]};
            assign {t0[13], t0[15]} = (in[13] > in[15]) ? {in[15], in[13]} : {in[13], in[15]};
            assign {t0[16], t0[18]} = (in[16] > in[18]) ? {in[18], in[16]} : {in[16], in[18]};
            assign {t0[17], t0[19]} = (in[17] > in[19]) ? {in[19], in[17]} : {in[17], in[19]};
            assign {t0[20], t0[22]} = (in[20] > in[22]) ? {in[22], in[20]} : {in[20], in[22]};
            assign {t0[21], t0[23]} = (in[21] > in[23]) ? {in[23], in[21]} : {in[21], in[23]};
            assign {t0[24], t0[26]} = (in[24] > in[26]) ? {in[26], in[24]} : {in[24], in[26]};
            assign {t0[25], t0[27]} = (in[25] > in[27]) ? {in[27], in[25]} : {in[25], in[27]};
            assign {t0[28], t0[30]} = (in[28] > in[30]) ? {in[30], in[28]} : {in[28], in[30]};
            assign {t0[29], t0[31]} = (in[29] > in[31]) ? {in[31], in[29]} : {in[29], in[31]};
            assign {t0[32], t0[34]} = (in[32] > in[34]) ? {in[34], in[32]} : {in[32], in[34]};
            assign {t0[33], t0[35]} = (in[33] > in[35]) ? {in[35], in[33]} : {in[33], in[35]};
            assign {t0[36], t0[38]} = (in[36] > in[38]) ? {in[38], in[36]} : {in[36], in[38]};
            assign {t0[37], t0[39]} = (in[37] > in[39]) ? {in[39], in[37]} : {in[37], in[39]};
            assign {t0[40], t0[42]} = (in[40] > in[42]) ? {in[42], in[40]} : {in[40], in[42]};
            assign {t0[41], t0[43]} = (in[41] > in[43]) ? {in[43], in[41]} : {in[41], in[43]};
            assign {t0[44], t0[46]} = (in[44] > in[46]) ? {in[46], in[44]} : {in[44], in[46]};
            assign {t0[45], t0[47]} = (in[45] > in[47]) ? {in[47], in[45]} : {in[45], in[47]};
            assign {t0[48], t0[50]} = (in[48] > in[50]) ? {in[50], in[48]} : {in[48], in[50]};
            assign {t0[49], t0[51]} = (in[49] > in[51]) ? {in[51], in[49]} : {in[49], in[51]};
            assign {t0[52], t0[54]} = (in[52] > in[54]) ? {in[54], in[52]} : {in[52], in[54]};
            assign {t0[53], t0[55]} = (in[53] > in[55]) ? {in[55], in[53]} : {in[53], in[55]};
            assign {t0[56], t0[58]} = (in[56] > in[58]) ? {in[58], in[56]} : {in[56], in[58]};
            assign {t0[57], t0[59]} = (in[57] > in[59]) ? {in[59], in[57]} : {in[57], in[59]};
            assign {t0[60], t0[62]} = (in[60] > in[62]) ? {in[62], in[60]} : {in[60], in[62]};
            assign {t0[61], t0[63]} = (in[61] > in[63]) ? {in[63], in[61]} : {in[61], in[63]};
            assign {t1[0], t1[1]} = (t0[0] > t0[1]) ? {t0[1], t0[0]} : {t0[0], t0[1]};
            assign {t1[2], t1[3]} = (t0[2] > t0[3]) ? {t0[3], t0[2]} : {t0[2], t0[3]};
            assign {t1[4], t1[5]} = (t0[4] > t0[5]) ? {t0[5], t0[4]} : {t0[4], t0[5]};
            assign {t1[6], t1[7]} = (t0[6] > t0[7]) ? {t0[7], t0[6]} : {t0[6], t0[7]};
            assign {t1[8], t1[9]} = (t0[8] > t0[9]) ? {t0[9], t0[8]} : {t0[8], t0[9]};
            assign {t1[10], t1[11]} = (t0[10] > t0[11]) ? {t0[11], t0[10]} : {t0[10], t0[11]};
            assign {t1[12], t1[13]} = (t0[12] > t0[13]) ? {t0[13], t0[12]} : {t0[12], t0[13]};
            assign {t1[14], t1[15]} = (t0[14] > t0[15]) ? {t0[15], t0[14]} : {t0[14], t0[15]};
            assign {t1[16], t1[17]} = (t0[16] > t0[17]) ? {t0[17], t0[16]} : {t0[16], t0[17]};
            assign {t1[18], t1[19]} = (t0[18] > t0[19]) ? {t0[19], t0[18]} : {t0[18], t0[19]};
            assign {t1[20], t1[21]} = (t0[20] > t0[21]) ? {t0[21], t0[20]} : {t0[20], t0[21]};
            assign {t1[22], t1[23]} = (t0[22] > t0[23]) ? {t0[23], t0[22]} : {t0[22], t0[23]};
            assign {t1[24], t1[25]} = (t0[24] > t0[25]) ? {t0[25], t0[24]} : {t0[24], t0[25]};
            assign {t1[26], t1[27]} = (t0[26] > t0[27]) ? {t0[27], t0[26]} : {t0[26], t0[27]};
            assign {t1[28], t1[29]} = (t0[28] > t0[29]) ? {t0[29], t0[28]} : {t0[28], t0[29]};
            assign {t1[30], t1[31]} = (t0[30] > t0[31]) ? {t0[31], t0[30]} : {t0[30], t0[31]};
            assign {t1[32], t1[33]} = (t0[32] > t0[33]) ? {t0[33], t0[32]} : {t0[32], t0[33]};
            assign {t1[34], t1[35]} = (t0[34] > t0[35]) ? {t0[35], t0[34]} : {t0[34], t0[35]};
            assign {t1[36], t1[37]} = (t0[36] > t0[37]) ? {t0[37], t0[36]} : {t0[36], t0[37]};
            assign {t1[38], t1[39]} = (t0[38] > t0[39]) ? {t0[39], t0[38]} : {t0[38], t0[39]};
            assign {t1[40], t1[41]} = (t0[40] > t0[41]) ? {t0[41], t0[40]} : {t0[40], t0[41]};
            assign {t1[42], t1[43]} = (t0[42] > t0[43]) ? {t0[43], t0[42]} : {t0[42], t0[43]};
            assign {t1[44], t1[45]} = (t0[44] > t0[45]) ? {t0[45], t0[44]} : {t0[44], t0[45]};
            assign {t1[46], t1[47]} = (t0[46] > t0[47]) ? {t0[47], t0[46]} : {t0[46], t0[47]};
            assign {t1[48], t1[49]} = (t0[48] > t0[49]) ? {t0[49], t0[48]} : {t0[48], t0[49]};
            assign {t1[50], t1[51]} = (t0[50] > t0[51]) ? {t0[51], t0[50]} : {t0[50], t0[51]};
            assign {t1[52], t1[53]} = (t0[52] > t0[53]) ? {t0[53], t0[52]} : {t0[52], t0[53]};
            assign {t1[54], t1[55]} = (t0[54] > t0[55]) ? {t0[55], t0[54]} : {t0[54], t0[55]};
            assign {t1[56], t1[57]} = (t0[56] > t0[57]) ? {t0[57], t0[56]} : {t0[56], t0[57]};
            assign {t1[58], t1[59]} = (t0[58] > t0[59]) ? {t0[59], t0[58]} : {t0[58], t0[59]};
            assign {t1[60], t1[61]} = (t0[60] > t0[61]) ? {t0[61], t0[60]} : {t0[60], t0[61]};
            assign {t1[62], t1[63]} = (t0[62] > t0[63]) ? {t0[63], t0[62]} : {t0[62], t0[63]};
            assign {t2[0], t2[20]} = (t1[0] > t1[20]) ? {t1[20], t1[0]} : {t1[0], t1[20]};
            assign {t2[1], t2[2]} = (t1[1] > t1[2]) ? {t1[2], t1[1]} : {t1[1], t1[2]};
            assign {t2[3], t2[23]} = (t1[3] > t1[23]) ? {t1[23], t1[3]} : {t1[3], t1[23]};
            assign {t2[4], t2[16]} = (t1[4] > t1[16]) ? {t1[16], t1[4]} : {t1[4], t1[16]};
            assign {t2[5], t2[6]} = (t1[5] > t1[6]) ? {t1[6], t1[5]} : {t1[5], t1[6]};
            assign {t2[7], t2[19]} = (t1[7] > t1[19]) ? {t1[19], t1[7]} : {t1[7], t1[19]};
            assign {t2[8], t2[48]} = (t1[8] > t1[48]) ? {t1[48], t1[8]} : {t1[8], t1[48]};
            assign {t2[9], t2[10]} = (t1[9] > t1[10]) ? {t1[10], t1[9]} : {t1[9], t1[10]};
            assign {t2[11], t2[51]} = (t1[11] > t1[51]) ? {t1[51], t1[11]} : {t1[11], t1[51]};
            assign {t2[12], t2[52]} = (t1[12] > t1[52]) ? {t1[52], t1[12]} : {t1[12], t1[52]};
            assign {t2[13], t2[14]} = (t1[13] > t1[14]) ? {t1[14], t1[13]} : {t1[13], t1[14]};
            assign {t2[15], t2[55]} = (t1[15] > t1[55]) ? {t1[55], t1[15]} : {t1[15], t1[55]};
            assign {t2[17], t2[18]} = (t1[17] > t1[18]) ? {t1[18], t1[17]} : {t1[17], t1[18]};
            assign {t2[21], t2[22]} = (t1[21] > t1[22]) ? {t1[22], t1[21]} : {t1[21], t1[22]};
            assign {t2[24], t2[28]} = (t1[24] > t1[28]) ? {t1[28], t1[24]} : {t1[24], t1[28]};
            assign {t2[25], t2[26]} = (t1[25] > t1[26]) ? {t1[26], t1[25]} : {t1[25], t1[26]};
            assign {t2[27], t2[31]} = (t1[27] > t1[31]) ? {t1[31], t1[27]} : {t1[27], t1[31]};
            assign {t2[29], t2[30]} = (t1[29] > t1[30]) ? {t1[30], t1[29]} : {t1[29], t1[30]};
            assign {t2[32], t2[36]} = (t1[32] > t1[36]) ? {t1[36], t1[32]} : {t1[32], t1[36]};
            assign {t2[33], t2[34]} = (t1[33] > t1[34]) ? {t1[34], t1[33]} : {t1[33], t1[34]};
            assign {t2[35], t2[39]} = (t1[35] > t1[39]) ? {t1[39], t1[35]} : {t1[35], t1[39]};
            assign {t2[37], t2[38]} = (t1[37] > t1[38]) ? {t1[38], t1[37]} : {t1[37], t1[38]};
            assign {t2[40], t2[60]} = (t1[40] > t1[60]) ? {t1[60], t1[40]} : {t1[40], t1[60]};
            assign {t2[41], t2[42]} = (t1[41] > t1[42]) ? {t1[42], t1[41]} : {t1[41], t1[42]};
            assign {t2[43], t2[63]} = (t1[43] > t1[63]) ? {t1[63], t1[43]} : {t1[43], t1[63]};
            assign {t2[44], t2[56]} = (t1[44] > t1[56]) ? {t1[56], t1[44]} : {t1[44], t1[56]};
            assign {t2[45], t2[46]} = (t1[45] > t1[46]) ? {t1[46], t1[45]} : {t1[45], t1[46]};
            assign {t2[47], t2[59]} = (t1[47] > t1[59]) ? {t1[59], t1[47]} : {t1[47], t1[59]};
            assign {t2[49], t2[50]} = (t1[49] > t1[50]) ? {t1[50], t1[49]} : {t1[49], t1[50]};
            assign {t2[53], t2[54]} = (t1[53] > t1[54]) ? {t1[54], t1[53]} : {t1[53], t1[54]};
            assign {t2[57], t2[58]} = (t1[57] > t1[58]) ? {t1[58], t1[57]} : {t1[57], t1[58]};
            assign {t2[61], t2[62]} = (t1[61] > t1[62]) ? {t1[62], t1[61]} : {t1[61], t1[62]};
            assign {t3[0], t3[8]} = (t2[0] > t2[8]) ? {t2[8], t2[0]} : {t2[0], t2[8]};
            assign {t3[1], t3[21]} = (t2[1] > t2[21]) ? {t2[21], t2[1]} : {t2[1], t2[21]};
            assign {t3[2], t3[22]} = (t2[2] > t2[22]) ? {t2[22], t2[2]} : {t2[2], t2[22]};
            assign {t3[3], t3[11]} = (t2[3] > t2[11]) ? {t2[11], t2[3]} : {t2[3], t2[11]};
            assign {t3[4], t3[40]} = (t2[4] > t2[40]) ? {t2[40], t2[4]} : {t2[4], t2[40]};
            assign {t3[5], t3[17]} = (t2[5] > t2[17]) ? {t2[17], t2[5]} : {t2[5], t2[17]};
            assign {t3[6], t3[18]} = (t2[6] > t2[18]) ? {t2[18], t2[6]} : {t2[6], t2[18]};
            assign {t3[7], t3[43]} = (t2[7] > t2[43]) ? {t2[43], t2[7]} : {t2[7], t2[43]};
            assign {t3[9], t3[49]} = (t2[9] > t2[49]) ? {t2[49], t2[9]} : {t2[9], t2[49]};
            assign {t3[10], t3[50]} = (t2[10] > t2[50]) ? {t2[50], t2[10]} : {t2[10], t2[50]};
            assign {t3[12], t3[24]} = (t2[12] > t2[24]) ? {t2[24], t2[12]} : {t2[12], t2[24]};
            assign {t3[13], t3[53]} = (t2[13] > t2[53]) ? {t2[53], t2[13]} : {t2[13], t2[53]};
            assign {t3[14], t3[54]} = (t2[14] > t2[54]) ? {t2[54], t2[14]} : {t2[14], t2[54]};
            assign {t3[15], t3[27]} = (t2[15] > t2[27]) ? {t2[27], t2[15]} : {t2[15], t2[27]};
            assign {t3[16], t3[28]} = (t2[16] > t2[28]) ? {t2[28], t2[16]} : {t2[16], t2[28]};
            assign {t3[19], t3[31]} = (t2[19] > t2[31]) ? {t2[31], t2[19]} : {t2[19], t2[31]};
            assign {t3[20], t3[56]} = (t2[20] > t2[56]) ? {t2[56], t2[20]} : {t2[20], t2[56]};
            assign {t3[23], t3[59]} = (t2[23] > t2[59]) ? {t2[59], t2[23]} : {t2[23], t2[59]};
            assign {t3[25], t3[29]} = (t2[25] > t2[29]) ? {t2[29], t2[25]} : {t2[25], t2[29]};
            assign {t3[26], t3[30]} = (t2[26] > t2[30]) ? {t2[30], t2[26]} : {t2[26], t2[30]};
            assign {t3[32], t3[44]} = (t2[32] > t2[44]) ? {t2[44], t2[32]} : {t2[32], t2[44]};
            assign {t3[33], t3[37]} = (t2[33] > t2[37]) ? {t2[37], t2[33]} : {t2[33], t2[37]};
            assign {t3[34], t3[38]} = (t2[34] > t2[38]) ? {t2[38], t2[34]} : {t2[34], t2[38]};
            assign {t3[35], t3[47]} = (t2[35] > t2[47]) ? {t2[47], t2[35]} : {t2[35], t2[47]};
            assign {t3[36], t3[48]} = (t2[36] > t2[48]) ? {t2[48], t2[36]} : {t2[36], t2[48]};
            assign {t3[39], t3[51]} = (t2[39] > t2[51]) ? {t2[51], t2[39]} : {t2[39], t2[51]};
            assign {t3[41], t3[61]} = (t2[41] > t2[61]) ? {t2[61], t2[41]} : {t2[41], t2[61]};
            assign {t3[42], t3[62]} = (t2[42] > t2[62]) ? {t2[62], t2[42]} : {t2[42], t2[62]};
            assign {t3[45], t3[57]} = (t2[45] > t2[57]) ? {t2[57], t2[45]} : {t2[45], t2[57]};
            assign {t3[46], t3[58]} = (t2[46] > t2[58]) ? {t2[58], t2[46]} : {t2[46], t2[58]};
            assign {t3[52], t3[60]} = (t2[52] > t2[60]) ? {t2[60], t2[52]} : {t2[52], t2[60]};
            assign {t3[55], t3[63]} = (t2[55] > t2[63]) ? {t2[63], t2[55]} : {t2[55], t2[63]};
            assign {t4[0], t4[32]} = (t3[0] > t3[32]) ? {t3[32], t3[0]} : {t3[0], t3[32]};
            assign {t4[1], t4[9]} = (t3[1] > t3[9]) ? {t3[9], t3[1]} : {t3[1], t3[9]};
            assign {t4[2], t4[10]} = (t3[2] > t3[10]) ? {t3[10], t3[2]} : {t3[2], t3[10]};
            assign {t4[3], t4[35]} = (t3[3] > t3[35]) ? {t3[35], t3[3]} : {t3[3], t3[35]};
            assign {t4[4], t4[12]} = (t3[4] > t3[12]) ? {t3[12], t3[4]} : {t3[4], t3[12]};
            assign {t4[5], t4[41]} = (t3[5] > t3[41]) ? {t3[41], t3[5]} : {t3[5], t3[41]};
            assign {t4[6], t4[42]} = (t3[6] > t3[42]) ? {t3[42], t3[6]} : {t3[6], t3[42]};
            assign {t4[7], t4[15]} = (t3[7] > t3[15]) ? {t3[15], t3[7]} : {t3[7], t3[15]};
            assign {t4[8], t4[44]} = (t3[8] > t3[44]) ? {t3[44], t3[8]} : {t3[8], t3[44]};
            assign {t4[11], t4[47]} = (t3[11] > t3[47]) ? {t3[47], t3[11]} : {t3[11], t3[47]};
            assign {t4[13], t4[25]} = (t3[13] > t3[25]) ? {t3[25], t3[13]} : {t3[13], t3[25]};
            assign {t4[14], t4[26]} = (t3[14] > t3[26]) ? {t3[26], t3[14]} : {t3[14], t3[26]};
            assign {t4[16], t4[52]} = (t3[16] > t3[52]) ? {t3[52], t3[16]} : {t3[16], t3[52]};
            assign {t4[17], t4[29]} = (t3[17] > t3[29]) ? {t3[29], t3[17]} : {t3[17], t3[29]};
            assign {t4[18], t4[30]} = (t3[18] > t3[30]) ? {t3[30], t3[18]} : {t3[18], t3[30]};
            assign {t4[19], t4[55]} = (t3[19] > t3[55]) ? {t3[55], t3[19]} : {t3[19], t3[55]};
            assign {t4[20], t4[36]} = (t3[20] > t3[36]) ? {t3[36], t3[20]} : {t3[20], t3[36]};
            assign {t4[21], t4[57]} = (t3[21] > t3[57]) ? {t3[57], t3[21]} : {t3[21], t3[57]};
            assign {t4[22], t4[58]} = (t3[22] > t3[58]) ? {t3[58], t3[22]} : {t3[22], t3[58]};
            assign {t4[23], t4[39]} = (t3[23] > t3[39]) ? {t3[39], t3[23]} : {t3[23], t3[39]};
            assign {t4[24], t4[40]} = (t3[24] > t3[40]) ? {t3[40], t3[24]} : {t3[24], t3[40]};
            assign {t4[27], t4[43]} = (t3[27] > t3[43]) ? {t3[43], t3[27]} : {t3[27], t3[43]};
            assign {t4[28], t4[60]} = (t3[28] > t3[60]) ? {t3[60], t3[28]} : {t3[28], t3[60]};
            assign {t4[31], t4[63]} = (t3[31] > t3[63]) ? {t3[63], t3[31]} : {t3[31], t3[63]};
            assign {t4[33], t4[45]} = (t3[33] > t3[45]) ? {t3[45], t3[33]} : {t3[33], t3[45]};
            assign {t4[34], t4[46]} = (t3[34] > t3[46]) ? {t3[46], t3[34]} : {t3[34], t3[46]};
            assign {t4[37], t4[49]} = (t3[37] > t3[49]) ? {t3[49], t3[37]} : {t3[37], t3[49]};
            assign {t4[38], t4[50]} = (t3[38] > t3[50]) ? {t3[50], t3[38]} : {t3[38], t3[50]};
            assign {t4[48], t4[56]} = (t3[48] > t3[56]) ? {t3[56], t3[48]} : {t3[48], t3[56]};
            assign {t4[51], t4[59]} = (t3[51] > t3[59]) ? {t3[59], t3[51]} : {t3[51], t3[59]};
            assign {t4[53], t4[61]} = (t3[53] > t3[61]) ? {t3[61], t3[53]} : {t3[53], t3[61]};
            assign {t4[54], t4[62]} = (t3[54] > t3[62]) ? {t3[62], t3[54]} : {t3[54], t3[62]};
            assign {t5[0], t5[4]} = (t4[0] > t4[4]) ? {t4[4], t4[0]} : {t4[0], t4[4]};
            assign {t5[1], t5[33]} = (t4[1] > t4[33]) ? {t4[33], t4[1]} : {t4[1], t4[33]};
            assign {t5[2], t5[34]} = (t4[2] > t4[34]) ? {t4[34], t4[2]} : {t4[2], t4[34]};
            assign {t5[3], t5[7]} = (t4[3] > t4[7]) ? {t4[7], t4[3]} : {t4[3], t4[7]};
            assign {t5[5], t5[13]} = (t4[5] > t4[13]) ? {t4[13], t4[5]} : {t4[5], t4[13]};
            assign {t5[6], t5[14]} = (t4[6] > t4[14]) ? {t4[14], t4[6]} : {t4[6], t4[14]};
            assign {t5[8], t5[16]} = (t4[8] > t4[16]) ? {t4[16], t4[8]} : {t4[8], t4[16]};
            assign {t5[9], t5[45]} = (t4[9] > t4[45]) ? {t4[45], t4[9]} : {t4[9], t4[45]};
            assign {t5[10], t5[46]} = (t4[10] > t4[46]) ? {t4[46], t4[10]} : {t4[10], t4[46]};
            assign {t5[11], t5[19]} = (t4[11] > t4[19]) ? {t4[19], t4[11]} : {t4[11], t4[19]};
            assign {t5[12], t5[32]} = (t4[12] > t4[32]) ? {t4[32], t4[12]} : {t4[12], t4[32]};
            assign {t5[15], t5[35]} = (t4[15] > t4[35]) ? {t4[35], t4[15]} : {t4[15], t4[35]};
            assign {t5[17], t5[53]} = (t4[17] > t4[53]) ? {t4[53], t4[17]} : {t4[17], t4[53]};
            assign {t5[18], t5[54]} = (t4[18] > t4[54]) ? {t4[54], t4[18]} : {t4[18], t4[54]};
            assign {t5[20], t5[24]} = (t4[20] > t4[24]) ? {t4[24], t4[20]} : {t4[20], t4[24]};
            assign {t5[21], t5[37]} = (t4[21] > t4[37]) ? {t4[37], t4[21]} : {t4[21], t4[37]};
            assign {t5[22], t5[38]} = (t4[22] > t4[38]) ? {t4[38], t4[22]} : {t4[22], t4[38]};
            assign {t5[23], t5[27]} = (t4[23] > t4[27]) ? {t4[27], t4[23]} : {t4[23], t4[27]};
            assign {t5[25], t5[41]} = (t4[25] > t4[41]) ? {t4[41], t4[25]} : {t4[25], t4[41]};
            assign {t5[26], t5[42]} = (t4[26] > t4[42]) ? {t4[42], t4[26]} : {t4[26], t4[42]};
            assign {t5[28], t5[48]} = (t4[28] > t4[48]) ? {t4[48], t4[28]} : {t4[28], t4[48]};
            assign {t5[29], t5[61]} = (t4[29] > t4[61]) ? {t4[61], t4[29]} : {t4[29], t4[61]};
            assign {t5[30], t5[62]} = (t4[30] > t4[62]) ? {t4[62], t4[30]} : {t4[30], t4[62]};
            assign {t5[31], t5[51]} = (t4[31] > t4[51]) ? {t4[51], t4[31]} : {t4[31], t4[51]};
            assign {t5[36], t5[40]} = (t4[36] > t4[40]) ? {t4[40], t4[36]} : {t4[36], t4[40]};
            assign {t5[39], t5[43]} = (t4[39] > t4[43]) ? {t4[43], t4[39]} : {t4[39], t4[43]};
            assign {t5[44], t5[52]} = (t4[44] > t4[52]) ? {t4[52], t4[44]} : {t4[44], t4[52]};
            assign {t5[47], t5[55]} = (t4[47] > t4[55]) ? {t4[55], t4[47]} : {t4[47], t4[55]};
            assign {t5[49], t5[57]} = (t4[49] > t4[57]) ? {t4[57], t4[49]} : {t4[49], t4[57]};
            assign {t5[50], t5[58]} = (t4[50] > t4[58]) ? {t4[58], t4[50]} : {t4[50], t4[58]};
            assign {t5[56], t5[60]} = (t4[56] > t4[60]) ? {t4[60], t4[56]} : {t4[56], t4[60]};
            assign {t5[59], t5[63]} = (t4[59] > t4[63]) ? {t4[63], t4[59]} : {t4[59], t4[63]};
            assign {t6[1], t6[5]} = (t5[1] > t5[5]) ? {t5[5], t5[1]} : {t5[1], t5[5]};
            assign {t6[2], t6[6]} = (t5[2] > t5[6]) ? {t5[6], t5[2]} : {t5[2], t5[6]};
            assign {t6[4], t6[12]} = (t5[4] > t5[12]) ? {t5[12], t5[4]} : {t5[4], t5[12]};
            assign {t6[7], t6[15]} = (t5[7] > t5[15]) ? {t5[15], t5[7]} : {t5[7], t5[15]};
            assign {t6[8], t6[20]} = (t5[8] > t5[20]) ? {t5[20], t5[8]} : {t5[8], t5[20]};
            assign {t6[9], t6[17]} = (t5[9] > t5[17]) ? {t5[17], t5[9]} : {t5[9], t5[17]};
            assign {t6[10], t6[18]} = (t5[10] > t5[18]) ? {t5[18], t5[10]} : {t5[10], t5[18]};
            assign {t6[11], t6[23]} = (t5[11] > t5[23]) ? {t5[23], t5[11]} : {t5[11], t5[23]};
            assign {t6[13], t6[33]} = (t5[13] > t5[33]) ? {t5[33], t5[13]} : {t5[13], t5[33]};
            assign {t6[14], t6[34]} = (t5[14] > t5[34]) ? {t5[34], t5[14]} : {t5[14], t5[34]};
            assign {t6[16], t6[32]} = (t5[16] > t5[32]) ? {t5[32], t5[16]} : {t5[16], t5[32]};
            assign {t6[19], t6[35]} = (t5[19] > t5[35]) ? {t5[35], t5[19]} : {t5[19], t5[35]};
            assign {t6[21], t6[25]} = (t5[21] > t5[25]) ? {t5[25], t5[21]} : {t5[21], t5[25]};
            assign {t6[22], t6[26]} = (t5[22] > t5[26]) ? {t5[26], t5[22]} : {t5[22], t5[26]};
            assign {t6[24], t6[36]} = (t5[24] > t5[36]) ? {t5[36], t5[24]} : {t5[24], t5[36]};
            assign {t6[27], t6[39]} = (t5[27] > t5[39]) ? {t5[39], t5[27]} : {t5[27], t5[39]};
            assign {t6[28], t6[44]} = (t5[28] > t5[44]) ? {t5[44], t5[28]} : {t5[28], t5[44]};
            assign {t6[29], t6[49]} = (t5[29] > t5[49]) ? {t5[49], t5[29]} : {t5[29], t5[49]};
            assign {t6[30], t6[50]} = (t5[30] > t5[50]) ? {t5[50], t5[30]} : {t5[30], t5[50]};
            assign {t6[31], t6[47]} = (t5[31] > t5[47]) ? {t5[47], t5[31]} : {t5[31], t5[47]};
            assign {t6[37], t6[41]} = (t5[37] > t5[41]) ? {t5[41], t5[37]} : {t5[37], t5[41]};
            assign {t6[38], t6[42]} = (t5[38] > t5[42]) ? {t5[42], t5[38]} : {t5[38], t5[42]};
            assign {t6[40], t6[52]} = (t5[40] > t5[52]) ? {t5[52], t5[40]} : {t5[40], t5[52]};
            assign {t6[43], t6[55]} = (t5[43] > t5[55]) ? {t5[55], t5[43]} : {t5[43], t5[55]};
            assign {t6[45], t6[53]} = (t5[45] > t5[53]) ? {t5[53], t5[45]} : {t5[45], t5[53]};
            assign {t6[46], t6[54]} = (t5[46] > t5[54]) ? {t5[54], t5[46]} : {t5[46], t5[54]};
            assign {t6[48], t6[56]} = (t5[48] > t5[56]) ? {t5[56], t5[48]} : {t5[48], t5[56]};
            assign {t6[51], t6[59]} = (t5[51] > t5[59]) ? {t5[59], t5[51]} : {t5[51], t5[59]};
            assign {t6[57], t6[61]} = (t5[57] > t5[61]) ? {t5[61], t5[57]} : {t5[57], t5[61]};
            assign {t6[58], t6[62]} = (t5[58] > t5[62]) ? {t5[62], t5[58]} : {t5[58], t5[62]};
            assign t6[0] = t5[0];
            assign t6[3] = t5[3];
            assign t6[60] = t5[60];
            assign t6[63] = t5[63];
            assign {t7[4], t7[8]} = (t6[4] > t6[8]) ? {t6[8], t6[4]} : {t6[4], t6[8]};
            assign {t7[5], t7[13]} = (t6[5] > t6[13]) ? {t6[13], t6[5]} : {t6[5], t6[13]};
            assign {t7[6], t7[14]} = (t6[6] > t6[14]) ? {t6[14], t6[6]} : {t6[6], t6[14]};
            assign {t7[7], t7[11]} = (t6[7] > t6[11]) ? {t6[11], t6[7]} : {t6[7], t6[11]};
            assign {t7[9], t7[21]} = (t6[9] > t6[21]) ? {t6[21], t6[9]} : {t6[9], t6[21]};
            assign {t7[10], t7[22]} = (t6[10] > t6[22]) ? {t6[22], t6[10]} : {t6[10], t6[22]};
            assign {t7[12], t7[20]} = (t6[12] > t6[20]) ? {t6[20], t6[12]} : {t6[12], t6[20]};
            assign {t7[15], t7[23]} = (t6[15] > t6[23]) ? {t6[23], t6[15]} : {t6[15], t6[23]};
            assign {t7[16], t7[44]} = (t6[16] > t6[44]) ? {t6[44], t6[16]} : {t6[16], t6[44]};
            assign {t7[17], t7[33]} = (t6[17] > t6[33]) ? {t6[33], t6[17]} : {t6[17], t6[33]};
            assign {t7[18], t7[34]} = (t6[18] > t6[34]) ? {t6[34], t6[18]} : {t6[18], t6[34]};
            assign {t7[19], t7[47]} = (t6[19] > t6[47]) ? {t6[47], t6[19]} : {t6[19], t6[47]};
            assign {t7[24], t7[32]} = (t6[24] > t6[32]) ? {t6[32], t6[24]} : {t6[24], t6[32]};
            assign {t7[25], t7[37]} = (t6[25] > t6[37]) ? {t6[37], t6[25]} : {t6[25], t6[37]};
            assign {t7[26], t7[38]} = (t6[26] > t6[38]) ? {t6[38], t6[26]} : {t6[26], t6[38]};
            assign {t7[27], t7[35]} = (t6[27] > t6[35]) ? {t6[35], t6[27]} : {t6[27], t6[35]};
            assign {t7[28], t7[36]} = (t6[28] > t6[36]) ? {t6[36], t6[28]} : {t6[28], t6[36]};
            assign {t7[29], t7[45]} = (t6[29] > t6[45]) ? {t6[45], t6[29]} : {t6[29], t6[45]};
            assign {t7[30], t7[46]} = (t6[30] > t6[46]) ? {t6[46], t6[30]} : {t6[30], t6[46]};
            assign {t7[31], t7[39]} = (t6[31] > t6[39]) ? {t6[39], t6[31]} : {t6[31], t6[39]};
            assign {t7[40], t7[48]} = (t6[40] > t6[48]) ? {t6[48], t6[40]} : {t6[40], t6[48]};
            assign {t7[41], t7[53]} = (t6[41] > t6[53]) ? {t6[53], t6[41]} : {t6[41], t6[53]};
            assign {t7[42], t7[54]} = (t6[42] > t6[54]) ? {t6[54], t6[42]} : {t6[42], t6[54]};
            assign {t7[43], t7[51]} = (t6[43] > t6[51]) ? {t6[51], t6[43]} : {t6[43], t6[51]};
            assign {t7[49], t7[57]} = (t6[49] > t6[57]) ? {t6[57], t6[49]} : {t6[49], t6[57]};
            assign {t7[50], t7[58]} = (t6[50] > t6[58]) ? {t6[58], t6[50]} : {t6[50], t6[58]};
            assign {t7[52], t7[56]} = (t6[52] > t6[56]) ? {t6[56], t6[52]} : {t6[52], t6[56]};
            assign {t7[55], t7[59]} = (t6[55] > t6[59]) ? {t6[59], t6[55]} : {t6[55], t6[59]};
            assign t7[0] = t6[0];
            assign t7[1] = t6[1];
            assign t7[2] = t6[2];
            assign t7[3] = t6[3];
            assign t7[60] = t6[60];
            assign t7[61] = t6[61];
            assign t7[62] = t6[62];
            assign t7[63] = t6[63];
            assign {t8[5], t8[9]} = (t7[5] > t7[9]) ? {t7[9], t7[5]} : {t7[5], t7[9]};
            assign {t8[6], t8[10]} = (t7[6] > t7[10]) ? {t7[10], t7[6]} : {t7[6], t7[10]};
            assign {t8[8], t8[12]} = (t7[8] > t7[12]) ? {t7[12], t7[8]} : {t7[8], t7[12]};
            assign {t8[11], t8[15]} = (t7[11] > t7[15]) ? {t7[15], t7[11]} : {t7[11], t7[15]};
            assign {t8[13], t8[21]} = (t7[13] > t7[21]) ? {t7[21], t7[13]} : {t7[13], t7[21]};
            assign {t8[14], t8[22]} = (t7[14] > t7[22]) ? {t7[22], t7[14]} : {t7[14], t7[22]};
            assign {t8[16], t8[20]} = (t7[16] > t7[20]) ? {t7[20], t7[16]} : {t7[16], t7[20]};
            assign {t8[17], t8[45]} = (t7[17] > t7[45]) ? {t7[45], t7[17]} : {t7[17], t7[45]};
            assign {t8[18], t8[46]} = (t7[18] > t7[46]) ? {t7[46], t7[18]} : {t7[18], t7[46]};
            assign {t8[19], t8[23]} = (t7[19] > t7[23]) ? {t7[23], t7[19]} : {t7[19], t7[23]};
            assign {t8[24], t8[28]} = (t7[24] > t7[28]) ? {t7[28], t7[24]} : {t7[24], t7[28]};
            assign {t8[25], t8[33]} = (t7[25] > t7[33]) ? {t7[33], t7[25]} : {t7[25], t7[33]};
            assign {t8[26], t8[34]} = (t7[26] > t7[34]) ? {t7[34], t7[26]} : {t7[26], t7[34]};
            assign {t8[27], t8[31]} = (t7[27] > t7[31]) ? {t7[31], t7[27]} : {t7[27], t7[31]};
            assign {t8[29], t8[37]} = (t7[29] > t7[37]) ? {t7[37], t7[29]} : {t7[29], t7[37]};
            assign {t8[30], t8[38]} = (t7[30] > t7[38]) ? {t7[38], t7[30]} : {t7[30], t7[38]};
            assign {t8[32], t8[36]} = (t7[32] > t7[36]) ? {t7[36], t7[32]} : {t7[32], t7[36]};
            assign {t8[35], t8[39]} = (t7[35] > t7[39]) ? {t7[39], t7[35]} : {t7[35], t7[39]};
            assign {t8[40], t8[44]} = (t7[40] > t7[44]) ? {t7[44], t7[40]} : {t7[40], t7[44]};
            assign {t8[41], t8[49]} = (t7[41] > t7[49]) ? {t7[49], t7[41]} : {t7[41], t7[49]};
            assign {t8[42], t8[50]} = (t7[42] > t7[50]) ? {t7[50], t7[42]} : {t7[42], t7[50]};
            assign {t8[43], t8[47]} = (t7[43] > t7[47]) ? {t7[47], t7[43]} : {t7[43], t7[47]};
            assign {t8[48], t8[52]} = (t7[48] > t7[52]) ? {t7[52], t7[48]} : {t7[48], t7[52]};
            assign {t8[51], t8[55]} = (t7[51] > t7[55]) ? {t7[55], t7[51]} : {t7[51], t7[55]};
            assign {t8[53], t8[57]} = (t7[53] > t7[57]) ? {t7[57], t7[53]} : {t7[53], t7[57]};
            assign {t8[54], t8[58]} = (t7[54] > t7[58]) ? {t7[58], t7[54]} : {t7[54], t7[58]};
            assign t8[0] = t7[0];
            assign t8[1] = t7[1];
            assign t8[2] = t7[2];
            assign t8[3] = t7[3];
            assign t8[4] = t7[4];
            assign t8[7] = t7[7];
            assign t8[56] = t7[56];
            assign t8[59] = t7[59];
            assign t8[60] = t7[60];
            assign t8[61] = t7[61];
            assign t8[62] = t7[62];
            assign t8[63] = t7[63];
            assign {t9[9], t9[13]} = (t8[9] > t8[13]) ? {t8[13], t8[9]} : {t8[9], t8[13]};
            assign {t9[10], t9[14]} = (t8[10] > t8[14]) ? {t8[14], t8[10]} : {t8[10], t8[14]};
            assign {t9[16], t9[24]} = (t8[16] > t8[24]) ? {t8[24], t8[16]} : {t8[16], t8[24]};
            assign {t9[17], t9[21]} = (t8[17] > t8[21]) ? {t8[21], t8[17]} : {t8[17], t8[21]};
            assign {t9[18], t9[22]} = (t8[18] > t8[22]) ? {t8[22], t8[18]} : {t8[18], t8[22]};
            assign {t9[19], t9[27]} = (t8[19] > t8[27]) ? {t8[27], t8[19]} : {t8[19], t8[27]};
            assign {t9[20], t9[28]} = (t8[20] > t8[28]) ? {t8[28], t8[20]} : {t8[20], t8[28]};
            assign {t9[23], t9[31]} = (t8[23] > t8[31]) ? {t8[31], t8[23]} : {t8[23], t8[31]};
            assign {t9[25], t9[29]} = (t8[25] > t8[29]) ? {t8[29], t8[25]} : {t8[25], t8[29]};
            assign {t9[26], t9[30]} = (t8[26] > t8[30]) ? {t8[30], t8[26]} : {t8[26], t8[30]};
            assign {t9[32], t9[40]} = (t8[32] > t8[40]) ? {t8[40], t8[32]} : {t8[32], t8[40]};
            assign {t9[33], t9[37]} = (t8[33] > t8[37]) ? {t8[37], t8[33]} : {t8[33], t8[37]};
            assign {t9[34], t9[38]} = (t8[34] > t8[38]) ? {t8[38], t8[34]} : {t8[34], t8[38]};
            assign {t9[35], t9[43]} = (t8[35] > t8[43]) ? {t8[43], t8[35]} : {t8[35], t8[43]};
            assign {t9[36], t9[44]} = (t8[36] > t8[44]) ? {t8[44], t8[36]} : {t8[36], t8[44]};
            assign {t9[39], t9[47]} = (t8[39] > t8[47]) ? {t8[47], t8[39]} : {t8[39], t8[47]};
            assign {t9[41], t9[45]} = (t8[41] > t8[45]) ? {t8[45], t8[41]} : {t8[41], t8[45]};
            assign {t9[42], t9[46]} = (t8[42] > t8[46]) ? {t8[46], t8[42]} : {t8[42], t8[46]};
            assign {t9[49], t9[53]} = (t8[49] > t8[53]) ? {t8[53], t8[49]} : {t8[49], t8[53]};
            assign {t9[50], t9[54]} = (t8[50] > t8[54]) ? {t8[54], t8[50]} : {t8[50], t8[54]};
            assign t9[0] = t8[0];
            assign t9[1] = t8[1];
            assign t9[2] = t8[2];
            assign t9[3] = t8[3];
            assign t9[4] = t8[4];
            assign t9[5] = t8[5];
            assign t9[6] = t8[6];
            assign t9[7] = t8[7];
            assign t9[8] = t8[8];
            assign t9[11] = t8[11];
            assign t9[12] = t8[12];
            assign t9[15] = t8[15];
            assign t9[48] = t8[48];
            assign t9[51] = t8[51];
            assign t9[52] = t8[52];
            assign t9[55] = t8[55];
            assign t9[56] = t8[56];
            assign t9[57] = t8[57];
            assign t9[58] = t8[58];
            assign t9[59] = t8[59];
            assign t9[60] = t8[60];
            assign t9[61] = t8[61];
            assign t9[62] = t8[62];
            assign t9[63] = t8[63];
            assign {t10[12], t10[16]} = (t9[12] > t9[16]) ? {t9[16], t9[12]} : {t9[12], t9[16]};
            assign {t10[15], t10[19]} = (t9[15] > t9[19]) ? {t9[19], t9[15]} : {t9[15], t9[19]};
            assign {t10[17], t10[25]} = (t9[17] > t9[25]) ? {t9[25], t9[17]} : {t9[17], t9[25]};
            assign {t10[18], t10[26]} = (t9[18] > t9[26]) ? {t9[26], t9[18]} : {t9[18], t9[26]};
            assign {t10[20], t10[24]} = (t9[20] > t9[24]) ? {t9[24], t9[20]} : {t9[20], t9[24]};
            assign {t10[21], t10[29]} = (t9[21] > t9[29]) ? {t9[29], t9[21]} : {t9[21], t9[29]};
            assign {t10[22], t10[30]} = (t9[22] > t9[30]) ? {t9[30], t9[22]} : {t9[22], t9[30]};
            assign {t10[23], t10[27]} = (t9[23] > t9[27]) ? {t9[27], t9[23]} : {t9[23], t9[27]};
            assign {t10[28], t10[32]} = (t9[28] > t9[32]) ? {t9[32], t9[28]} : {t9[28], t9[32]};
            assign {t10[31], t10[35]} = (t9[31] > t9[35]) ? {t9[35], t9[31]} : {t9[31], t9[35]};
            assign {t10[33], t10[41]} = (t9[33] > t9[41]) ? {t9[41], t9[33]} : {t9[33], t9[41]};
            assign {t10[34], t10[42]} = (t9[34] > t9[42]) ? {t9[42], t9[34]} : {t9[34], t9[42]};
            assign {t10[36], t10[40]} = (t9[36] > t9[40]) ? {t9[40], t9[36]} : {t9[36], t9[40]};
            assign {t10[37], t10[45]} = (t9[37] > t9[45]) ? {t9[45], t9[37]} : {t9[37], t9[45]};
            assign {t10[38], t10[46]} = (t9[38] > t9[46]) ? {t9[46], t9[38]} : {t9[38], t9[46]};
            assign {t10[39], t10[43]} = (t9[39] > t9[43]) ? {t9[43], t9[39]} : {t9[39], t9[43]};
            assign {t10[44], t10[48]} = (t9[44] > t9[48]) ? {t9[48], t9[44]} : {t9[44], t9[48]};
            assign {t10[47], t10[51]} = (t9[47] > t9[51]) ? {t9[51], t9[47]} : {t9[47], t9[51]};
            assign t10[0] = t9[0];
            assign t10[1] = t9[1];
            assign t10[2] = t9[2];
            assign t10[3] = t9[3];
            assign t10[4] = t9[4];
            assign t10[5] = t9[5];
            assign t10[6] = t9[6];
            assign t10[7] = t9[7];
            assign t10[8] = t9[8];
            assign t10[9] = t9[9];
            assign t10[10] = t9[10];
            assign t10[11] = t9[11];
            assign t10[13] = t9[13];
            assign t10[14] = t9[14];
            assign t10[49] = t9[49];
            assign t10[50] = t9[50];
            assign t10[52] = t9[52];
            assign t10[53] = t9[53];
            assign t10[54] = t9[54];
            assign t10[55] = t9[55];
            assign t10[56] = t9[56];
            assign t10[57] = t9[57];
            assign t10[58] = t9[58];
            assign t10[59] = t9[59];
            assign t10[60] = t9[60];
            assign t10[61] = t9[61];
            assign t10[62] = t9[62];
            assign t10[63] = t9[63];
            assign {t11[1], t11[16]} = (t10[1] > t10[16]) ? {t10[16], t10[1]} : {t10[1], t10[16]};
            assign {t11[2], t11[32]} = (t10[2] > t10[32]) ? {t10[32], t10[2]} : {t10[2], t10[32]};
            assign {t11[5], t11[20]} = (t10[5] > t10[20]) ? {t10[20], t10[5]} : {t10[5], t10[20]};
            assign {t11[6], t11[36]} = (t10[6] > t10[36]) ? {t10[36], t10[6]} : {t10[6], t10[36]};
            assign {t11[9], t11[24]} = (t10[9] > t10[24]) ? {t10[24], t10[9]} : {t10[9], t10[24]};
            assign {t11[10], t11[40]} = (t10[10] > t10[40]) ? {t10[40], t10[10]} : {t10[10], t10[40]};
            assign {t11[13], t11[17]} = (t10[13] > t10[17]) ? {t10[17], t10[13]} : {t10[13], t10[17]};
            assign {t11[14], t11[18]} = (t10[14] > t10[18]) ? {t10[18], t10[14]} : {t10[14], t10[18]};
            assign {t11[21], t11[25]} = (t10[21] > t10[25]) ? {t10[25], t10[21]} : {t10[21], t10[25]};
            assign {t11[22], t11[26]} = (t10[22] > t10[26]) ? {t10[26], t10[22]} : {t10[22], t10[26]};
            assign {t11[23], t11[53]} = (t10[23] > t10[53]) ? {t10[53], t10[23]} : {t10[23], t10[53]};
            assign {t11[27], t11[57]} = (t10[27] > t10[57]) ? {t10[57], t10[27]} : {t10[27], t10[57]};
            assign {t11[29], t11[33]} = (t10[29] > t10[33]) ? {t10[33], t10[29]} : {t10[29], t10[33]};
            assign {t11[30], t11[34]} = (t10[30] > t10[34]) ? {t10[34], t10[30]} : {t10[30], t10[34]};
            assign {t11[31], t11[61]} = (t10[31] > t10[61]) ? {t10[61], t10[31]} : {t10[31], t10[61]};
            assign {t11[37], t11[41]} = (t10[37] > t10[41]) ? {t10[41], t10[37]} : {t10[37], t10[41]};
            assign {t11[38], t11[42]} = (t10[38] > t10[42]) ? {t10[42], t10[38]} : {t10[38], t10[42]};
            assign {t11[39], t11[54]} = (t10[39] > t10[54]) ? {t10[54], t10[39]} : {t10[39], t10[54]};
            assign {t11[43], t11[58]} = (t10[43] > t10[58]) ? {t10[58], t10[43]} : {t10[43], t10[58]};
            assign {t11[45], t11[49]} = (t10[45] > t10[49]) ? {t10[49], t10[45]} : {t10[45], t10[49]};
            assign {t11[46], t11[50]} = (t10[46] > t10[50]) ? {t10[50], t10[46]} : {t10[46], t10[50]};
            assign {t11[47], t11[62]} = (t10[47] > t10[62]) ? {t10[62], t10[47]} : {t10[47], t10[62]};
            assign t11[0] = t10[0];
            assign t11[3] = t10[3];
            assign t11[4] = t10[4];
            assign t11[7] = t10[7];
            assign t11[8] = t10[8];
            assign t11[11] = t10[11];
            assign t11[12] = t10[12];
            assign t11[15] = t10[15];
            assign t11[19] = t10[19];
            assign t11[28] = t10[28];
            assign t11[35] = t10[35];
            assign t11[44] = t10[44];
            assign t11[48] = t10[48];
            assign t11[51] = t10[51];
            assign t11[52] = t10[52];
            assign t11[55] = t10[55];
            assign t11[56] = t10[56];
            assign t11[59] = t10[59];
            assign t11[60] = t10[60];
            assign t11[63] = t10[63];
            assign {t12[1], t12[4]} = (t11[1] > t11[4]) ? {t11[4], t11[1]} : {t11[1], t11[4]};
            assign {t12[2], t12[8]} = (t11[2] > t11[8]) ? {t11[8], t11[2]} : {t11[2], t11[8]};
            assign {t12[3], t12[33]} = (t11[3] > t11[33]) ? {t11[33], t11[3]} : {t11[3], t11[33]};
            assign {t12[6], t12[12]} = (t11[6] > t11[12]) ? {t11[12], t11[6]} : {t11[6], t11[12]};
            assign {t12[7], t12[37]} = (t11[7] > t11[37]) ? {t11[37], t11[7]} : {t11[7], t11[37]};
            assign {t12[10], t12[24]} = (t11[10] > t11[24]) ? {t11[24], t11[10]} : {t11[10], t11[24]};
            assign {t12[11], t12[41]} = (t11[11] > t11[41]) ? {t11[41], t11[11]} : {t11[11], t11[41]};
            assign {t12[13], t12[28]} = (t11[13] > t11[28]) ? {t11[28], t11[13]} : {t11[13], t11[28]};
            assign {t12[14], t12[44]} = (t11[14] > t11[44]) ? {t11[44], t11[14]} : {t11[14], t11[44]};
            assign {t12[15], t12[45]} = (t11[15] > t11[45]) ? {t11[45], t11[15]} : {t11[15], t11[45]};
            assign {t12[18], t12[48]} = (t11[18] > t11[48]) ? {t11[48], t11[18]} : {t11[18], t11[48]};
            assign {t12[19], t12[49]} = (t11[19] > t11[49]) ? {t11[49], t11[19]} : {t11[19], t11[49]};
            assign {t12[21], t12[36]} = (t11[21] > t11[36]) ? {t11[36], t11[21]} : {t11[21], t11[36]};
            assign {t12[22], t12[52]} = (t11[22] > t11[52]) ? {t11[52], t11[22]} : {t11[22], t11[52]};
            assign {t12[26], t12[56]} = (t11[26] > t11[56]) ? {t11[56], t11[26]} : {t11[26], t11[56]};
            assign {t12[27], t12[42]} = (t11[27] > t11[42]) ? {t11[42], t11[27]} : {t11[27], t11[42]};
            assign {t12[30], t12[60]} = (t11[30] > t11[60]) ? {t11[60], t11[30]} : {t11[30], t11[60]};
            assign {t12[35], t12[50]} = (t11[35] > t11[50]) ? {t11[50], t11[35]} : {t11[35], t11[50]};
            assign {t12[39], t12[53]} = (t11[39] > t11[53]) ? {t11[53], t11[39]} : {t11[39], t11[53]};
            assign {t12[51], t12[57]} = (t11[51] > t11[57]) ? {t11[57], t11[51]} : {t11[51], t11[57]};
            assign {t12[55], t12[61]} = (t11[55] > t11[61]) ? {t11[61], t11[55]} : {t11[55], t11[61]};
            assign {t12[59], t12[62]} = (t11[59] > t11[62]) ? {t11[62], t11[59]} : {t11[59], t11[62]};
            assign t12[0] = t11[0];
            assign t12[5] = t11[5];
            assign t12[9] = t11[9];
            assign t12[16] = t11[16];
            assign t12[17] = t11[17];
            assign t12[20] = t11[20];
            assign t12[23] = t11[23];
            assign t12[25] = t11[25];
            assign t12[29] = t11[29];
            assign t12[31] = t11[31];
            assign t12[32] = t11[32];
            assign t12[34] = t11[34];
            assign t12[38] = t11[38];
            assign t12[40] = t11[40];
            assign t12[43] = t11[43];
            assign t12[46] = t11[46];
            assign t12[47] = t11[47];
            assign t12[54] = t11[54];
            assign t12[58] = t11[58];
            assign t12[63] = t11[63];
            assign {t13[2], t13[4]} = (t12[2] > t12[4]) ? {t12[4], t12[2]} : {t12[2], t12[4]};
            assign {t13[3], t13[17]} = (t12[3] > t12[17]) ? {t12[17], t12[3]} : {t12[3], t12[17]};
            assign {t13[5], t13[6]} = (t12[5] > t12[6]) ? {t12[6], t12[5]} : {t12[5], t12[6]};
            assign {t13[7], t13[22]} = (t12[7] > t12[22]) ? {t12[22], t12[7]} : {t12[7], t12[22]};
            assign {t13[8], t13[16]} = (t12[8] > t12[16]) ? {t12[16], t12[8]} : {t12[8], t12[16]};
            assign {t13[11], t13[25]} = (t12[11] > t12[25]) ? {t12[25], t12[11]} : {t12[11], t12[25]};
            assign {t13[12], t13[20]} = (t12[12] > t12[20]) ? {t12[20], t12[12]} : {t12[12], t12[20]};
            assign {t13[14], t13[28]} = (t12[14] > t12[28]) ? {t12[28], t12[14]} : {t12[14], t12[28]};
            assign {t13[15], t13[29]} = (t12[15] > t12[29]) ? {t12[29], t12[15]} : {t12[15], t12[29]};
            assign {t13[18], t13[32]} = (t12[18] > t12[32]) ? {t12[32], t12[18]} : {t12[18], t12[32]};
            assign {t13[19], t13[33]} = (t12[19] > t12[33]) ? {t12[33], t12[19]} : {t12[19], t12[33]};
            assign {t13[23], t13[37]} = (t12[23] > t12[37]) ? {t12[37], t12[23]} : {t12[23], t12[37]};
            assign {t13[26], t13[40]} = (t12[26] > t12[40]) ? {t12[40], t12[26]} : {t12[26], t12[40]};
            assign {t13[30], t13[44]} = (t12[30] > t12[44]) ? {t12[44], t12[30]} : {t12[30], t12[44]};
            assign {t13[31], t13[45]} = (t12[31] > t12[45]) ? {t12[45], t12[31]} : {t12[31], t12[45]};
            assign {t13[34], t13[48]} = (t12[34] > t12[48]) ? {t12[48], t12[34]} : {t12[34], t12[48]};
            assign {t13[35], t13[49]} = (t12[35] > t12[49]) ? {t12[49], t12[35]} : {t12[35], t12[49]};
            assign {t13[38], t13[52]} = (t12[38] > t12[52]) ? {t12[52], t12[38]} : {t12[38], t12[52]};
            assign {t13[41], t13[56]} = (t12[41] > t12[56]) ? {t12[56], t12[41]} : {t12[41], t12[56]};
            assign {t13[43], t13[51]} = (t12[43] > t12[51]) ? {t12[51], t12[43]} : {t12[43], t12[51]};
            assign {t13[46], t13[60]} = (t12[46] > t12[60]) ? {t12[60], t12[46]} : {t12[46], t12[60]};
            assign {t13[47], t13[55]} = (t12[47] > t12[55]) ? {t12[55], t12[47]} : {t12[47], t12[55]};
            assign {t13[57], t13[58]} = (t12[57] > t12[58]) ? {t12[58], t12[57]} : {t12[57], t12[58]};
            assign {t13[59], t13[61]} = (t12[59] > t12[61]) ? {t12[61], t12[59]} : {t12[59], t12[61]};
            assign t13[0] = t12[0];
            assign t13[1] = t12[1];
            assign t13[9] = t12[9];
            assign t13[10] = t12[10];
            assign t13[13] = t12[13];
            assign t13[21] = t12[21];
            assign t13[24] = t12[24];
            assign t13[27] = t12[27];
            assign t13[36] = t12[36];
            assign t13[39] = t12[39];
            assign t13[42] = t12[42];
            assign t13[50] = t12[50];
            assign t13[53] = t12[53];
            assign t13[54] = t12[54];
            assign t13[62] = t12[62];
            assign t13[63] = t12[63];
            assign {t14[3], t14[18]} = (t13[3] > t13[18]) ? {t13[18], t13[3]} : {t13[3], t13[18]};
            assign {t14[7], t14[21]} = (t13[7] > t13[21]) ? {t13[21], t13[7]} : {t13[7], t13[21]};
            assign {t14[11], t14[32]} = (t13[11] > t13[32]) ? {t13[32], t13[11]} : {t13[11], t13[32]};
            assign {t14[15], t14[30]} = (t13[15] > t13[30]) ? {t13[30], t13[15]} : {t13[15], t13[30]};
            assign {t14[17], t14[26]} = (t13[17] > t13[26]) ? {t13[26], t13[17]} : {t13[17], t13[26]};
            assign {t14[19], t14[25]} = (t13[19] > t13[25]) ? {t13[25], t13[19]} : {t13[19], t13[25]};
            assign {t14[22], t14[36]} = (t13[22] > t13[36]) ? {t13[36], t13[22]} : {t13[22], t13[36]};
            assign {t14[23], t14[29]} = (t13[23] > t13[29]) ? {t13[29], t13[23]} : {t13[23], t13[29]};
            assign {t14[27], t14[41]} = (t13[27] > t13[41]) ? {t13[41], t13[27]} : {t13[27], t13[41]};
            assign {t14[31], t14[52]} = (t13[31] > t13[52]) ? {t13[52], t13[31]} : {t13[31], t13[52]};
            assign {t14[33], t14[48]} = (t13[33] > t13[48]) ? {t13[48], t13[33]} : {t13[33], t13[48]};
            assign {t14[34], t14[40]} = (t13[34] > t13[40]) ? {t13[40], t13[34]} : {t13[34], t13[40]};
            assign {t14[37], t14[46]} = (t13[37] > t13[46]) ? {t13[46], t13[37]} : {t13[37], t13[46]};
            assign {t14[38], t14[44]} = (t13[38] > t13[44]) ? {t13[44], t13[38]} : {t13[38], t13[44]};
            assign {t14[42], t14[56]} = (t13[42] > t13[56]) ? {t13[56], t13[42]} : {t13[42], t13[56]};
            assign {t14[45], t14[60]} = (t13[45] > t13[60]) ? {t13[60], t13[45]} : {t13[45], t13[60]};
            assign t14[0] = t13[0];
            assign t14[1] = t13[1];
            assign t14[2] = t13[2];
            assign t14[4] = t13[4];
            assign t14[5] = t13[5];
            assign t14[6] = t13[6];
            assign t14[8] = t13[8];
            assign t14[9] = t13[9];
            assign t14[10] = t13[10];
            assign t14[12] = t13[12];
            assign t14[13] = t13[13];
            assign t14[14] = t13[14];
            assign t14[16] = t13[16];
            assign t14[20] = t13[20];
            assign t14[24] = t13[24];
            assign t14[28] = t13[28];
            assign t14[35] = t13[35];
            assign t14[39] = t13[39];
            assign t14[43] = t13[43];
            assign t14[47] = t13[47];
            assign t14[49] = t13[49];
            assign t14[50] = t13[50];
            assign t14[51] = t13[51];
            assign t14[53] = t13[53];
            assign t14[54] = t13[54];
            assign t14[55] = t13[55];
            assign t14[57] = t13[57];
            assign t14[58] = t13[58];
            assign t14[59] = t13[59];
            assign t14[61] = t13[61];
            assign t14[62] = t13[62];
            assign t14[63] = t13[63];
            assign {t15[3], t15[16]} = (t14[3] > t14[16]) ? {t14[16], t14[3]} : {t14[3], t14[16]};
            assign {t15[7], t15[20]} = (t14[7] > t14[20]) ? {t14[20], t14[7]} : {t14[7], t14[20]};
            assign {t15[11], t15[24]} = (t14[11] > t14[24]) ? {t14[24], t14[11]} : {t14[11], t14[24]};
            assign {t15[15], t15[21]} = (t14[15] > t14[21]) ? {t14[21], t14[15]} : {t14[15], t14[21]};
            assign {t15[17], t15[18]} = (t14[17] > t14[18]) ? {t14[18], t14[17]} : {t14[17], t14[18]};
            assign {t15[19], t15[34]} = (t14[19] > t14[34]) ? {t14[34], t14[19]} : {t14[19], t14[34]};
            assign {t15[22], t15[28]} = (t14[22] > t14[28]) ? {t14[28], t14[22]} : {t14[22], t14[28]};
            assign {t15[23], t15[38]} = (t14[23] > t14[38]) ? {t14[38], t14[23]} : {t14[23], t14[38]};
            assign {t15[25], t15[40]} = (t14[25] > t14[40]) ? {t14[40], t14[25]} : {t14[25], t14[40]};
            assign {t15[26], t15[32]} = (t14[26] > t14[32]) ? {t14[32], t14[26]} : {t14[26], t14[32]};
            assign {t15[27], t15[33]} = (t14[27] > t14[33]) ? {t14[33], t14[27]} : {t14[27], t14[33]};
            assign {t15[29], t15[44]} = (t14[29] > t14[44]) ? {t14[44], t14[29]} : {t14[29], t14[44]};
            assign {t15[30], t15[36]} = (t14[30] > t14[36]) ? {t14[36], t14[30]} : {t14[30], t14[36]};
            assign {t15[31], t15[37]} = (t14[31] > t14[37]) ? {t14[37], t14[31]} : {t14[31], t14[37]};
            assign {t15[35], t15[41]} = (t14[35] > t14[41]) ? {t14[41], t14[35]} : {t14[35], t14[41]};
            assign {t15[39], t15[52]} = (t14[39] > t14[52]) ? {t14[52], t14[39]} : {t14[39], t14[52]};
            assign {t15[42], t15[48]} = (t14[42] > t14[48]) ? {t14[48], t14[42]} : {t14[42], t14[48]};
            assign {t15[43], t15[56]} = (t14[43] > t14[56]) ? {t14[56], t14[43]} : {t14[43], t14[56]};
            assign {t15[45], t15[46]} = (t14[45] > t14[46]) ? {t14[46], t14[45]} : {t14[45], t14[46]};
            assign {t15[47], t15[60]} = (t14[47] > t14[60]) ? {t14[60], t14[47]} : {t14[47], t14[60]};
            assign t15[0] = t14[0];
            assign t15[1] = t14[1];
            assign t15[2] = t14[2];
            assign t15[4] = t14[4];
            assign t15[5] = t14[5];
            assign t15[6] = t14[6];
            assign t15[8] = t14[8];
            assign t15[9] = t14[9];
            assign t15[10] = t14[10];
            assign t15[12] = t14[12];
            assign t15[13] = t14[13];
            assign t15[14] = t14[14];
            assign t15[49] = t14[49];
            assign t15[50] = t14[50];
            assign t15[51] = t14[51];
            assign t15[53] = t14[53];
            assign t15[54] = t14[54];
            assign t15[55] = t14[55];
            assign t15[57] = t14[57];
            assign t15[58] = t14[58];
            assign t15[59] = t14[59];
            assign t15[61] = t14[61];
            assign t15[62] = t14[62];
            assign t15[63] = t14[63];
            assign {t16[3], t16[9]} = (t15[3] > t15[9]) ? {t15[9], t15[3]} : {t15[3], t15[9]};
            assign {t16[7], t16[13]} = (t15[7] > t15[13]) ? {t15[13], t15[7]} : {t15[7], t15[13]};
            assign {t16[10], t16[16]} = (t15[10] > t15[16]) ? {t15[16], t15[10]} : {t15[10], t15[16]};
            assign {t16[11], t16[17]} = (t15[11] > t15[17]) ? {t15[17], t15[11]} : {t15[11], t15[17]};
            assign {t16[14], t16[20]} = (t15[14] > t15[20]) ? {t15[20], t15[14]} : {t15[14], t15[20]};
            assign {t16[15], t16[22]} = (t15[15] > t15[22]) ? {t15[22], t15[15]} : {t15[15], t15[22]};
            assign {t16[18], t16[24]} = (t15[18] > t15[24]) ? {t15[24], t15[18]} : {t15[18], t15[24]};
            assign {t16[19], t16[26]} = (t15[19] > t15[26]) ? {t15[26], t15[19]} : {t15[19], t15[26]};
            assign {t16[21], t16[28]} = (t15[21] > t15[28]) ? {t15[28], t15[21]} : {t15[21], t15[28]};
            assign {t16[23], t16[30]} = (t15[23] > t15[30]) ? {t15[30], t15[23]} : {t15[23], t15[30]};
            assign {t16[25], t16[32]} = (t15[25] > t15[32]) ? {t15[32], t15[25]} : {t15[25], t15[32]};
            assign {t16[27], t16[34]} = (t15[27] > t15[34]) ? {t15[34], t15[27]} : {t15[27], t15[34]};
            assign {t16[29], t16[36]} = (t15[29] > t15[36]) ? {t15[36], t15[29]} : {t15[29], t15[36]};
            assign {t16[31], t16[38]} = (t15[31] > t15[38]) ? {t15[38], t15[31]} : {t15[31], t15[38]};
            assign {t16[33], t16[40]} = (t15[33] > t15[40]) ? {t15[40], t15[33]} : {t15[33], t15[40]};
            assign {t16[35], t16[42]} = (t15[35] > t15[42]) ? {t15[42], t15[35]} : {t15[35], t15[42]};
            assign {t16[37], t16[44]} = (t15[37] > t15[44]) ? {t15[44], t15[37]} : {t15[37], t15[44]};
            assign {t16[39], t16[45]} = (t15[39] > t15[45]) ? {t15[45], t15[39]} : {t15[39], t15[45]};
            assign {t16[41], t16[48]} = (t15[41] > t15[48]) ? {t15[48], t15[41]} : {t15[41], t15[48]};
            assign {t16[43], t16[49]} = (t15[43] > t15[49]) ? {t15[49], t15[43]} : {t15[43], t15[49]};
            assign {t16[46], t16[52]} = (t15[46] > t15[52]) ? {t15[52], t15[46]} : {t15[46], t15[52]};
            assign {t16[47], t16[53]} = (t15[47] > t15[53]) ? {t15[53], t15[47]} : {t15[47], t15[53]};
            assign {t16[50], t16[56]} = (t15[50] > t15[56]) ? {t15[56], t15[50]} : {t15[50], t15[56]};
            assign {t16[54], t16[60]} = (t15[54] > t15[60]) ? {t15[60], t15[54]} : {t15[54], t15[60]};
            assign t16[0] = t15[0];
            assign t16[1] = t15[1];
            assign t16[2] = t15[2];
            assign t16[4] = t15[4];
            assign t16[5] = t15[5];
            assign t16[6] = t15[6];
            assign t16[8] = t15[8];
            assign t16[12] = t15[12];
            assign t16[51] = t15[51];
            assign t16[55] = t15[55];
            assign t16[57] = t15[57];
            assign t16[58] = t15[58];
            assign t16[59] = t15[59];
            assign t16[61] = t15[61];
            assign t16[62] = t15[62];
            assign t16[63] = t15[63];
            assign {t17[3], t17[8]} = (t16[3] > t16[8]) ? {t16[8], t16[3]} : {t16[3], t16[8]};
            assign {t17[7], t17[10]} = (t16[7] > t16[10]) ? {t16[10], t16[7]} : {t16[7], t16[10]};
            assign {t17[9], t17[12]} = (t16[9] > t16[12]) ? {t16[12], t16[9]} : {t16[9], t16[12]};
            assign {t17[11], t17[16]} = (t16[11] > t16[16]) ? {t16[16], t16[11]} : {t16[11], t16[16]};
            assign {t17[13], t17[14]} = (t16[13] > t16[14]) ? {t16[14], t16[13]} : {t16[13], t16[14]};
            assign {t17[15], t17[17]} = (t16[15] > t16[17]) ? {t16[17], t16[15]} : {t16[15], t16[17]};
            assign {t17[18], t17[20]} = (t16[18] > t16[20]) ? {t16[20], t16[18]} : {t16[18], t16[20]};
            assign {t17[19], t17[22]} = (t16[19] > t16[22]) ? {t16[22], t16[19]} : {t16[19], t16[22]};
            assign {t17[21], t17[24]} = (t16[21] > t16[24]) ? {t16[24], t16[21]} : {t16[21], t16[24]};
            assign {t17[23], t17[26]} = (t16[23] > t16[26]) ? {t16[26], t16[23]} : {t16[23], t16[26]};
            assign {t17[25], t17[28]} = (t16[25] > t16[28]) ? {t16[28], t16[25]} : {t16[25], t16[28]};
            assign {t17[27], t17[29]} = (t16[27] > t16[29]) ? {t16[29], t16[27]} : {t16[27], t16[29]};
            assign {t17[30], t17[32]} = (t16[30] > t16[32]) ? {t16[32], t16[30]} : {t16[30], t16[32]};
            assign {t17[31], t17[33]} = (t16[31] > t16[33]) ? {t16[33], t16[31]} : {t16[31], t16[33]};
            assign {t17[34], t17[36]} = (t16[34] > t16[36]) ? {t16[36], t16[34]} : {t16[34], t16[36]};
            assign {t17[35], t17[38]} = (t16[35] > t16[38]) ? {t16[38], t16[35]} : {t16[35], t16[38]};
            assign {t17[37], t17[40]} = (t16[37] > t16[40]) ? {t16[40], t16[37]} : {t16[37], t16[40]};
            assign {t17[39], t17[42]} = (t16[39] > t16[42]) ? {t16[42], t16[39]} : {t16[39], t16[42]};
            assign {t17[41], t17[44]} = (t16[41] > t16[44]) ? {t16[44], t16[41]} : {t16[41], t16[44]};
            assign {t17[43], t17[45]} = (t16[43] > t16[45]) ? {t16[45], t16[43]} : {t16[43], t16[45]};
            assign {t17[46], t17[48]} = (t16[46] > t16[48]) ? {t16[48], t16[46]} : {t16[46], t16[48]};
            assign {t17[47], t17[52]} = (t16[47] > t16[52]) ? {t16[52], t16[47]} : {t16[47], t16[52]};
            assign {t17[49], t17[50]} = (t16[49] > t16[50]) ? {t16[50], t16[49]} : {t16[49], t16[50]};
            assign {t17[51], t17[54]} = (t16[51] > t16[54]) ? {t16[54], t16[51]} : {t16[51], t16[54]};
            assign {t17[53], t17[56]} = (t16[53] > t16[56]) ? {t16[56], t16[53]} : {t16[53], t16[56]};
            assign {t17[55], t17[60]} = (t16[55] > t16[60]) ? {t16[60], t16[55]} : {t16[55], t16[60]};
            assign t17[0] = t16[0];
            assign t17[1] = t16[1];
            assign t17[2] = t16[2];
            assign t17[4] = t16[4];
            assign t17[5] = t16[5];
            assign t17[6] = t16[6];
            assign t17[57] = t16[57];
            assign t17[58] = t16[58];
            assign t17[59] = t16[59];
            assign t17[61] = t16[61];
            assign t17[62] = t16[62];
            assign t17[63] = t16[63];
            assign {t18[3], t18[5]} = (t17[3] > t17[5]) ? {t17[5], t17[3]} : {t17[3], t17[5]};
            assign {t18[6], t18[8]} = (t17[6] > t17[8]) ? {t17[8], t17[6]} : {t17[6], t17[8]};
            assign {t18[7], t18[9]} = (t17[7] > t17[9]) ? {t17[9], t17[7]} : {t17[7], t17[9]};
            assign {t18[10], t18[12]} = (t17[10] > t17[12]) ? {t17[12], t17[10]} : {t17[10], t17[12]};
            assign {t18[11], t18[13]} = (t17[11] > t17[13]) ? {t17[13], t17[11]} : {t17[11], t17[13]};
            assign {t18[14], t18[16]} = (t17[14] > t17[16]) ? {t17[16], t17[14]} : {t17[14], t17[16]};
            assign {t18[15], t18[18]} = (t17[15] > t17[18]) ? {t17[18], t17[15]} : {t17[15], t17[18]};
            assign {t18[17], t18[20]} = (t17[17] > t17[20]) ? {t17[20], t17[17]} : {t17[17], t17[20]};
            assign {t18[19], t18[21]} = (t17[19] > t17[21]) ? {t17[21], t17[19]} : {t17[19], t17[21]};
            assign {t18[22], t18[24]} = (t17[22] > t17[24]) ? {t17[24], t17[22]} : {t17[22], t17[24]};
            assign {t18[23], t18[25]} = (t17[23] > t17[25]) ? {t17[25], t17[23]} : {t17[23], t17[25]};
            assign {t18[26], t18[28]} = (t17[26] > t17[28]) ? {t17[28], t17[26]} : {t17[26], t17[28]};
            assign {t18[27], t18[30]} = (t17[27] > t17[30]) ? {t17[30], t17[27]} : {t17[27], t17[30]};
            assign {t18[29], t18[32]} = (t17[29] > t17[32]) ? {t17[32], t17[29]} : {t17[29], t17[32]};
            assign {t18[31], t18[34]} = (t17[31] > t17[34]) ? {t17[34], t17[31]} : {t17[31], t17[34]};
            assign {t18[33], t18[36]} = (t17[33] > t17[36]) ? {t17[36], t17[33]} : {t17[33], t17[36]};
            assign {t18[35], t18[37]} = (t17[35] > t17[37]) ? {t17[37], t17[35]} : {t17[35], t17[37]};
            assign {t18[38], t18[40]} = (t17[38] > t17[40]) ? {t17[40], t17[38]} : {t17[38], t17[40]};
            assign {t18[39], t18[41]} = (t17[39] > t17[41]) ? {t17[41], t17[39]} : {t17[39], t17[41]};
            assign {t18[42], t18[44]} = (t17[42] > t17[44]) ? {t17[44], t17[42]} : {t17[42], t17[44]};
            assign {t18[43], t18[46]} = (t17[43] > t17[46]) ? {t17[46], t17[43]} : {t17[43], t17[46]};
            assign {t18[45], t18[48]} = (t17[45] > t17[48]) ? {t17[48], t17[45]} : {t17[45], t17[48]};
            assign {t18[47], t18[49]} = (t17[47] > t17[49]) ? {t17[49], t17[47]} : {t17[47], t17[49]};
            assign {t18[50], t18[52]} = (t17[50] > t17[52]) ? {t17[52], t17[50]} : {t17[50], t17[52]};
            assign {t18[51], t18[53]} = (t17[51] > t17[53]) ? {t17[53], t17[51]} : {t17[51], t17[53]};
            assign {t18[54], t18[56]} = (t17[54] > t17[56]) ? {t17[56], t17[54]} : {t17[54], t17[56]};
            assign {t18[55], t18[57]} = (t17[55] > t17[57]) ? {t17[57], t17[55]} : {t17[55], t17[57]};
            assign {t18[58], t18[60]} = (t17[58] > t17[60]) ? {t17[60], t17[58]} : {t17[58], t17[60]};
            assign t18[0] = t17[0];
            assign t18[1] = t17[1];
            assign t18[2] = t17[2];
            assign t18[4] = t17[4];
            assign t18[59] = t17[59];
            assign t18[61] = t17[61];
            assign t18[62] = t17[62];
            assign t18[63] = t17[63];
            assign {t19[3], t19[4]} = (t18[3] > t18[4]) ? {t18[4], t18[3]} : {t18[3], t18[4]};
            assign {t19[5], t19[6]} = (t18[5] > t18[6]) ? {t18[6], t18[5]} : {t18[5], t18[6]};
            assign {t19[7], t19[8]} = (t18[7] > t18[8]) ? {t18[8], t18[7]} : {t18[7], t18[8]};
            assign {t19[9], t19[10]} = (t18[9] > t18[10]) ? {t18[10], t18[9]} : {t18[9], t18[10]};
            assign {t19[11], t19[12]} = (t18[11] > t18[12]) ? {t18[12], t18[11]} : {t18[11], t18[12]};
            assign {t19[13], t19[14]} = (t18[13] > t18[14]) ? {t18[14], t18[13]} : {t18[13], t18[14]};
            assign {t19[15], t19[16]} = (t18[15] > t18[16]) ? {t18[16], t18[15]} : {t18[15], t18[16]};
            assign {t19[17], t19[18]} = (t18[17] > t18[18]) ? {t18[18], t18[17]} : {t18[17], t18[18]};
            assign {t19[19], t19[20]} = (t18[19] > t18[20]) ? {t18[20], t18[19]} : {t18[19], t18[20]};
            assign {t19[21], t19[22]} = (t18[21] > t18[22]) ? {t18[22], t18[21]} : {t18[21], t18[22]};
            assign {t19[23], t19[24]} = (t18[23] > t18[24]) ? {t18[24], t18[23]} : {t18[23], t18[24]};
            assign {t19[25], t19[26]} = (t18[25] > t18[26]) ? {t18[26], t18[25]} : {t18[25], t18[26]};
            assign {t19[27], t19[28]} = (t18[27] > t18[28]) ? {t18[28], t18[27]} : {t18[27], t18[28]};
            assign {t19[29], t19[30]} = (t18[29] > t18[30]) ? {t18[30], t18[29]} : {t18[29], t18[30]};
            assign {t19[31], t19[32]} = (t18[31] > t18[32]) ? {t18[32], t18[31]} : {t18[31], t18[32]};
            assign {t19[33], t19[34]} = (t18[33] > t18[34]) ? {t18[34], t18[33]} : {t18[33], t18[34]};
            assign {t19[35], t19[36]} = (t18[35] > t18[36]) ? {t18[36], t18[35]} : {t18[35], t18[36]};
            assign {t19[37], t19[38]} = (t18[37] > t18[38]) ? {t18[38], t18[37]} : {t18[37], t18[38]};
            assign {t19[39], t19[40]} = (t18[39] > t18[40]) ? {t18[40], t18[39]} : {t18[39], t18[40]};
            assign {t19[41], t19[42]} = (t18[41] > t18[42]) ? {t18[42], t18[41]} : {t18[41], t18[42]};
            assign {t19[43], t19[44]} = (t18[43] > t18[44]) ? {t18[44], t18[43]} : {t18[43], t18[44]};
            assign {t19[45], t19[46]} = (t18[45] > t18[46]) ? {t18[46], t18[45]} : {t18[45], t18[46]};
            assign {t19[47], t19[48]} = (t18[47] > t18[48]) ? {t18[48], t18[47]} : {t18[47], t18[48]};
            assign {t19[49], t19[50]} = (t18[49] > t18[50]) ? {t18[50], t18[49]} : {t18[49], t18[50]};
            assign {t19[51], t19[52]} = (t18[51] > t18[52]) ? {t18[52], t18[51]} : {t18[51], t18[52]};
            assign {t19[53], t19[54]} = (t18[53] > t18[54]) ? {t18[54], t18[53]} : {t18[53], t18[54]};
            assign {t19[55], t19[56]} = (t18[55] > t18[56]) ? {t18[56], t18[55]} : {t18[55], t18[56]};
            assign {t19[57], t19[58]} = (t18[57] > t18[58]) ? {t18[58], t18[57]} : {t18[57], t18[58]};
            assign {t19[59], t19[60]} = (t18[59] > t18[60]) ? {t18[60], t18[59]} : {t18[59], t18[60]};
            assign t19[0] = t18[0];
            assign t19[1] = t18[1];
            assign t19[2] = t18[2];
            assign t19[61] = t18[61];
            assign t19[62] = t18[62];
            assign t19[63] = t18[63];

            if (DIRECTION == 0) begin
                always_ff @( posedge clk ) begin
                    out <= t19;
                end 
            end else begin
                for (i = 0; i < SIZE; i++) begin
                    always_ff @ ( posedge clk ) begin
                        out[i] <= t19[SIZE-i-1];
                    end
                end
            end
        end
    endgenerate
endmodule